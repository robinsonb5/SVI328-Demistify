
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"e0",x"80",x"00",x"00"),
     1 => (x"00",x"00",x"00",x"60"),
     2 => (x"08",x"08",x"08",x"00"),
     3 => (x"00",x"08",x"08",x"08"),
     4 => (x"60",x"00",x"00",x"00"),
     5 => (x"00",x"00",x"00",x"60"),
     6 => (x"18",x"30",x"60",x"40"),
     7 => (x"01",x"03",x"06",x"0c"),
     8 => (x"59",x"7f",x"3e",x"00"),
     9 => (x"00",x"3e",x"7f",x"4d"),
    10 => (x"7f",x"06",x"04",x"00"),
    11 => (x"00",x"00",x"00",x"7f"),
    12 => (x"71",x"63",x"42",x"00"),
    13 => (x"00",x"46",x"4f",x"59"),
    14 => (x"49",x"63",x"22",x"00"),
    15 => (x"00",x"36",x"7f",x"49"),
    16 => (x"13",x"16",x"1c",x"18"),
    17 => (x"00",x"10",x"7f",x"7f"),
    18 => (x"45",x"67",x"27",x"00"),
    19 => (x"00",x"39",x"7d",x"45"),
    20 => (x"4b",x"7e",x"3c",x"00"),
    21 => (x"00",x"30",x"79",x"49"),
    22 => (x"71",x"01",x"01",x"00"),
    23 => (x"00",x"07",x"0f",x"79"),
    24 => (x"49",x"7f",x"36",x"00"),
    25 => (x"00",x"36",x"7f",x"49"),
    26 => (x"49",x"4f",x"06",x"00"),
    27 => (x"00",x"1e",x"3f",x"69"),
    28 => (x"66",x"00",x"00",x"00"),
    29 => (x"00",x"00",x"00",x"66"),
    30 => (x"e6",x"80",x"00",x"00"),
    31 => (x"00",x"00",x"00",x"66"),
    32 => (x"14",x"08",x"08",x"00"),
    33 => (x"00",x"22",x"22",x"14"),
    34 => (x"14",x"14",x"14",x"00"),
    35 => (x"00",x"14",x"14",x"14"),
    36 => (x"14",x"22",x"22",x"00"),
    37 => (x"00",x"08",x"08",x"14"),
    38 => (x"51",x"03",x"02",x"00"),
    39 => (x"00",x"06",x"0f",x"59"),
    40 => (x"5d",x"41",x"7f",x"3e"),
    41 => (x"00",x"1e",x"1f",x"55"),
    42 => (x"09",x"7f",x"7e",x"00"),
    43 => (x"00",x"7e",x"7f",x"09"),
    44 => (x"49",x"7f",x"7f",x"00"),
    45 => (x"00",x"36",x"7f",x"49"),
    46 => (x"63",x"3e",x"1c",x"00"),
    47 => (x"00",x"41",x"41",x"41"),
    48 => (x"41",x"7f",x"7f",x"00"),
    49 => (x"00",x"1c",x"3e",x"63"),
    50 => (x"49",x"7f",x"7f",x"00"),
    51 => (x"00",x"41",x"41",x"49"),
    52 => (x"09",x"7f",x"7f",x"00"),
    53 => (x"00",x"01",x"01",x"09"),
    54 => (x"41",x"7f",x"3e",x"00"),
    55 => (x"00",x"7a",x"7b",x"49"),
    56 => (x"08",x"7f",x"7f",x"00"),
    57 => (x"00",x"7f",x"7f",x"08"),
    58 => (x"7f",x"41",x"00",x"00"),
    59 => (x"00",x"00",x"41",x"7f"),
    60 => (x"40",x"60",x"20",x"00"),
    61 => (x"00",x"3f",x"7f",x"40"),
    62 => (x"1c",x"08",x"7f",x"7f"),
    63 => (x"00",x"41",x"63",x"36"),
    64 => (x"40",x"7f",x"7f",x"00"),
    65 => (x"00",x"40",x"40",x"40"),
    66 => (x"0c",x"06",x"7f",x"7f"),
    67 => (x"00",x"7f",x"7f",x"06"),
    68 => (x"0c",x"06",x"7f",x"7f"),
    69 => (x"00",x"7f",x"7f",x"18"),
    70 => (x"41",x"7f",x"3e",x"00"),
    71 => (x"00",x"3e",x"7f",x"41"),
    72 => (x"09",x"7f",x"7f",x"00"),
    73 => (x"00",x"06",x"0f",x"09"),
    74 => (x"61",x"41",x"7f",x"3e"),
    75 => (x"00",x"40",x"7e",x"7f"),
    76 => (x"09",x"7f",x"7f",x"00"),
    77 => (x"00",x"66",x"7f",x"19"),
    78 => (x"4d",x"6f",x"26",x"00"),
    79 => (x"00",x"32",x"7b",x"59"),
    80 => (x"7f",x"01",x"01",x"00"),
    81 => (x"00",x"01",x"01",x"7f"),
    82 => (x"40",x"7f",x"3f",x"00"),
    83 => (x"00",x"3f",x"7f",x"40"),
    84 => (x"70",x"3f",x"0f",x"00"),
    85 => (x"00",x"0f",x"3f",x"70"),
    86 => (x"18",x"30",x"7f",x"7f"),
    87 => (x"00",x"7f",x"7f",x"30"),
    88 => (x"1c",x"36",x"63",x"41"),
    89 => (x"41",x"63",x"36",x"1c"),
    90 => (x"7c",x"06",x"03",x"01"),
    91 => (x"01",x"03",x"06",x"7c"),
    92 => (x"4d",x"59",x"71",x"61"),
    93 => (x"00",x"41",x"43",x"47"),
    94 => (x"7f",x"7f",x"00",x"00"),
    95 => (x"00",x"00",x"41",x"41"),
    96 => (x"0c",x"06",x"03",x"01"),
    97 => (x"40",x"60",x"30",x"18"),
    98 => (x"41",x"41",x"00",x"00"),
    99 => (x"00",x"00",x"7f",x"7f"),
   100 => (x"03",x"06",x"0c",x"08"),
   101 => (x"00",x"08",x"0c",x"06"),
   102 => (x"80",x"80",x"80",x"80"),
   103 => (x"00",x"80",x"80",x"80"),
   104 => (x"03",x"00",x"00",x"00"),
   105 => (x"00",x"00",x"04",x"07"),
   106 => (x"54",x"74",x"20",x"00"),
   107 => (x"00",x"78",x"7c",x"54"),
   108 => (x"44",x"7f",x"7f",x"00"),
   109 => (x"00",x"38",x"7c",x"44"),
   110 => (x"44",x"7c",x"38",x"00"),
   111 => (x"00",x"00",x"44",x"44"),
   112 => (x"44",x"7c",x"38",x"00"),
   113 => (x"00",x"7f",x"7f",x"44"),
   114 => (x"54",x"7c",x"38",x"00"),
   115 => (x"00",x"18",x"5c",x"54"),
   116 => (x"7f",x"7e",x"04",x"00"),
   117 => (x"00",x"00",x"05",x"05"),
   118 => (x"a4",x"bc",x"18",x"00"),
   119 => (x"00",x"7c",x"fc",x"a4"),
   120 => (x"04",x"7f",x"7f",x"00"),
   121 => (x"00",x"78",x"7c",x"04"),
   122 => (x"3d",x"00",x"00",x"00"),
   123 => (x"00",x"00",x"40",x"7d"),
   124 => (x"80",x"80",x"80",x"00"),
   125 => (x"00",x"00",x"7d",x"fd"),
   126 => (x"10",x"7f",x"7f",x"00"),
   127 => (x"00",x"44",x"6c",x"38"),
   128 => (x"3f",x"00",x"00",x"00"),
   129 => (x"00",x"00",x"40",x"7f"),
   130 => (x"18",x"0c",x"7c",x"7c"),
   131 => (x"00",x"78",x"7c",x"0c"),
   132 => (x"04",x"7c",x"7c",x"00"),
   133 => (x"00",x"78",x"7c",x"04"),
   134 => (x"44",x"7c",x"38",x"00"),
   135 => (x"00",x"38",x"7c",x"44"),
   136 => (x"24",x"fc",x"fc",x"00"),
   137 => (x"00",x"18",x"3c",x"24"),
   138 => (x"24",x"3c",x"18",x"00"),
   139 => (x"00",x"fc",x"fc",x"24"),
   140 => (x"04",x"7c",x"7c",x"00"),
   141 => (x"00",x"08",x"0c",x"04"),
   142 => (x"54",x"5c",x"48",x"00"),
   143 => (x"00",x"20",x"74",x"54"),
   144 => (x"7f",x"3f",x"04",x"00"),
   145 => (x"00",x"00",x"44",x"44"),
   146 => (x"40",x"7c",x"3c",x"00"),
   147 => (x"00",x"7c",x"7c",x"40"),
   148 => (x"60",x"3c",x"1c",x"00"),
   149 => (x"00",x"1c",x"3c",x"60"),
   150 => (x"30",x"60",x"7c",x"3c"),
   151 => (x"00",x"3c",x"7c",x"60"),
   152 => (x"10",x"38",x"6c",x"44"),
   153 => (x"00",x"44",x"6c",x"38"),
   154 => (x"e0",x"bc",x"1c",x"00"),
   155 => (x"00",x"1c",x"3c",x"60"),
   156 => (x"74",x"64",x"44",x"00"),
   157 => (x"00",x"44",x"4c",x"5c"),
   158 => (x"3e",x"08",x"08",x"00"),
   159 => (x"00",x"41",x"41",x"77"),
   160 => (x"7f",x"00",x"00",x"00"),
   161 => (x"00",x"00",x"00",x"7f"),
   162 => (x"77",x"41",x"41",x"00"),
   163 => (x"00",x"08",x"08",x"3e"),
   164 => (x"03",x"01",x"01",x"02"),
   165 => (x"00",x"01",x"02",x"02"),
   166 => (x"7f",x"7f",x"7f",x"7f"),
   167 => (x"00",x"7f",x"7f",x"7f"),
   168 => (x"1c",x"1c",x"08",x"08"),
   169 => (x"7f",x"7f",x"3e",x"3e"),
   170 => (x"3e",x"3e",x"7f",x"7f"),
   171 => (x"08",x"08",x"1c",x"1c"),
   172 => (x"7c",x"18",x"10",x"00"),
   173 => (x"00",x"10",x"18",x"7c"),
   174 => (x"7c",x"30",x"10",x"00"),
   175 => (x"00",x"10",x"30",x"7c"),
   176 => (x"60",x"60",x"30",x"10"),
   177 => (x"00",x"06",x"1e",x"78"),
   178 => (x"18",x"3c",x"66",x"42"),
   179 => (x"00",x"42",x"66",x"3c"),
   180 => (x"c2",x"6a",x"38",x"78"),
   181 => (x"00",x"38",x"6c",x"c6"),
   182 => (x"60",x"00",x"00",x"60"),
   183 => (x"00",x"60",x"00",x"00"),
   184 => (x"5c",x"5b",x"5e",x"0e"),
   185 => (x"86",x"fc",x"0e",x"5d"),
   186 => (x"f7",x"c2",x"7e",x"71"),
   187 => (x"c0",x"4c",x"bf",x"e0"),
   188 => (x"c4",x"1e",x"c0",x"4b"),
   189 => (x"c4",x"02",x"ab",x"66"),
   190 => (x"c2",x"4d",x"c0",x"87"),
   191 => (x"75",x"4d",x"c1",x"87"),
   192 => (x"ee",x"49",x"73",x"1e"),
   193 => (x"86",x"c8",x"87",x"e3"),
   194 => (x"ef",x"49",x"e0",x"c0"),
   195 => (x"a4",x"c4",x"87",x"ec"),
   196 => (x"f0",x"49",x"6a",x"4a"),
   197 => (x"ca",x"f1",x"87",x"f3"),
   198 => (x"c1",x"84",x"cc",x"87"),
   199 => (x"ab",x"b7",x"c8",x"83"),
   200 => (x"87",x"cd",x"ff",x"04"),
   201 => (x"4d",x"26",x"8e",x"fc"),
   202 => (x"4b",x"26",x"4c",x"26"),
   203 => (x"71",x"1e",x"4f",x"26"),
   204 => (x"e4",x"f7",x"c2",x"4a"),
   205 => (x"e4",x"f7",x"c2",x"5a"),
   206 => (x"49",x"78",x"c7",x"48"),
   207 => (x"26",x"87",x"e1",x"fe"),
   208 => (x"1e",x"73",x"1e",x"4f"),
   209 => (x"0b",x"fc",x"4b",x"71"),
   210 => (x"4a",x"73",x"0b",x"7b"),
   211 => (x"c0",x"c1",x"9a",x"c1"),
   212 => (x"c7",x"ed",x"49",x"a2"),
   213 => (x"d8",x"da",x"c2",x"87"),
   214 => (x"26",x"4b",x"26",x"5b"),
   215 => (x"4a",x"71",x"1e",x"4f"),
   216 => (x"72",x"1e",x"66",x"c4"),
   217 => (x"87",x"fb",x"eb",x"49"),
   218 => (x"4f",x"26",x"8e",x"fc"),
   219 => (x"48",x"d4",x"ff",x"1e"),
   220 => (x"ff",x"78",x"ff",x"c3"),
   221 => (x"e1",x"c0",x"48",x"d0"),
   222 => (x"48",x"d4",x"ff",x"78"),
   223 => (x"48",x"71",x"78",x"c1"),
   224 => (x"d4",x"ff",x"30",x"c4"),
   225 => (x"d0",x"ff",x"78",x"08"),
   226 => (x"78",x"e0",x"c0",x"48"),
   227 => (x"5e",x"0e",x"4f",x"26"),
   228 => (x"0e",x"5d",x"5c",x"5b"),
   229 => (x"7e",x"c0",x"86",x"f4"),
   230 => (x"ec",x"48",x"a6",x"c8"),
   231 => (x"80",x"fc",x"78",x"bf"),
   232 => (x"bf",x"e0",x"f7",x"c2"),
   233 => (x"e8",x"f7",x"c2",x"78"),
   234 => (x"bf",x"e8",x"4c",x"bf"),
   235 => (x"d4",x"da",x"c2",x"4d"),
   236 => (x"f9",x"e3",x"49",x"bf"),
   237 => (x"e8",x"49",x"c7",x"87"),
   238 => (x"49",x"70",x"87",x"f1"),
   239 => (x"d0",x"05",x"99",x"c2"),
   240 => (x"cc",x"da",x"c2",x"87"),
   241 => (x"b9",x"ff",x"49",x"bf"),
   242 => (x"c1",x"99",x"66",x"c8"),
   243 => (x"f9",x"c1",x"02",x"99"),
   244 => (x"49",x"e8",x"cf",x"87"),
   245 => (x"70",x"87",x"c1",x"cb"),
   246 => (x"e8",x"49",x"c7",x"4b"),
   247 => (x"98",x"70",x"87",x"cd"),
   248 => (x"c8",x"87",x"c9",x"05"),
   249 => (x"99",x"c1",x"49",x"66"),
   250 => (x"87",x"fe",x"c0",x"02"),
   251 => (x"ec",x"48",x"a6",x"c8"),
   252 => (x"f9",x"e2",x"78",x"bf"),
   253 => (x"ca",x"49",x"73",x"87"),
   254 => (x"98",x"70",x"87",x"ea"),
   255 => (x"c2",x"87",x"d7",x"02"),
   256 => (x"49",x"bf",x"c8",x"da"),
   257 => (x"da",x"c2",x"b9",x"c1"),
   258 => (x"fd",x"71",x"59",x"cc"),
   259 => (x"e8",x"cf",x"87",x"de"),
   260 => (x"87",x"c4",x"ca",x"49"),
   261 => (x"49",x"c7",x"4b",x"70"),
   262 => (x"70",x"87",x"d0",x"e7"),
   263 => (x"cb",x"ff",x"05",x"98"),
   264 => (x"49",x"66",x"c8",x"87"),
   265 => (x"ff",x"05",x"99",x"c1"),
   266 => (x"da",x"c2",x"87",x"c2"),
   267 => (x"c1",x"4a",x"bf",x"d4"),
   268 => (x"d8",x"da",x"c2",x"ba"),
   269 => (x"7a",x"0a",x"fc",x"5a"),
   270 => (x"c1",x"9a",x"c1",x"0a"),
   271 => (x"e9",x"49",x"a2",x"c0"),
   272 => (x"da",x"c1",x"87",x"da"),
   273 => (x"87",x"e3",x"e6",x"49"),
   274 => (x"da",x"c2",x"7e",x"c1"),
   275 => (x"66",x"c8",x"48",x"cc"),
   276 => (x"d4",x"da",x"c2",x"78"),
   277 => (x"e9",x"c0",x"05",x"bf"),
   278 => (x"c3",x"49",x"75",x"87"),
   279 => (x"1e",x"71",x"99",x"ff"),
   280 => (x"f8",x"fb",x"49",x"c0"),
   281 => (x"c8",x"49",x"75",x"87"),
   282 => (x"1e",x"71",x"29",x"b7"),
   283 => (x"ec",x"fb",x"49",x"c1"),
   284 => (x"c3",x"86",x"c8",x"87"),
   285 => (x"f2",x"e5",x"49",x"fd"),
   286 => (x"49",x"fa",x"c3",x"87"),
   287 => (x"c7",x"87",x"ec",x"e5"),
   288 => (x"49",x"75",x"87",x"f5"),
   289 => (x"c8",x"99",x"ff",x"c3"),
   290 => (x"b5",x"71",x"2d",x"b7"),
   291 => (x"c0",x"02",x"9d",x"75"),
   292 => (x"a6",x"c8",x"87",x"e4"),
   293 => (x"bf",x"c8",x"ff",x"48"),
   294 => (x"49",x"66",x"c8",x"78"),
   295 => (x"bf",x"d0",x"da",x"c2"),
   296 => (x"a9",x"e0",x"c2",x"89"),
   297 => (x"87",x"c4",x"c0",x"03"),
   298 => (x"87",x"d0",x"4d",x"c0"),
   299 => (x"48",x"d0",x"da",x"c2"),
   300 => (x"c0",x"78",x"66",x"c8"),
   301 => (x"da",x"c2",x"87",x"c6"),
   302 => (x"78",x"c0",x"48",x"d0"),
   303 => (x"99",x"c8",x"49",x"75"),
   304 => (x"87",x"ce",x"c0",x"05"),
   305 => (x"e4",x"49",x"f5",x"c3"),
   306 => (x"49",x"70",x"87",x"e1"),
   307 => (x"c0",x"02",x"99",x"c2"),
   308 => (x"f7",x"c2",x"87",x"e7"),
   309 => (x"c0",x"02",x"bf",x"e4"),
   310 => (x"c1",x"48",x"87",x"ca"),
   311 => (x"e8",x"f7",x"c2",x"88"),
   312 => (x"87",x"d3",x"c0",x"58"),
   313 => (x"c1",x"48",x"66",x"c4"),
   314 => (x"7e",x"70",x"80",x"e0"),
   315 => (x"c0",x"02",x"bf",x"6e"),
   316 => (x"ff",x"4b",x"87",x"c5"),
   317 => (x"c1",x"0f",x"73",x"49"),
   318 => (x"c4",x"49",x"75",x"7e"),
   319 => (x"ce",x"c0",x"05",x"99"),
   320 => (x"49",x"f2",x"c3",x"87"),
   321 => (x"70",x"87",x"e4",x"e3"),
   322 => (x"02",x"99",x"c2",x"49"),
   323 => (x"c2",x"87",x"eb",x"c0"),
   324 => (x"7e",x"bf",x"e4",x"f7"),
   325 => (x"b7",x"c7",x"48",x"6e"),
   326 => (x"cb",x"c0",x"03",x"a8"),
   327 => (x"c1",x"48",x"6e",x"87"),
   328 => (x"e8",x"f7",x"c2",x"80"),
   329 => (x"87",x"d0",x"c0",x"58"),
   330 => (x"c1",x"4a",x"66",x"c4"),
   331 => (x"02",x"6a",x"82",x"e0"),
   332 => (x"4b",x"87",x"c5",x"c0"),
   333 => (x"0f",x"73",x"49",x"fe"),
   334 => (x"fd",x"c3",x"7e",x"c1"),
   335 => (x"87",x"eb",x"e2",x"49"),
   336 => (x"99",x"c2",x"49",x"70"),
   337 => (x"87",x"e6",x"c0",x"02"),
   338 => (x"bf",x"e4",x"f7",x"c2"),
   339 => (x"87",x"c9",x"c0",x"02"),
   340 => (x"48",x"e4",x"f7",x"c2"),
   341 => (x"d3",x"c0",x"78",x"c0"),
   342 => (x"48",x"66",x"c4",x"87"),
   343 => (x"70",x"80",x"e0",x"c1"),
   344 => (x"02",x"bf",x"6e",x"7e"),
   345 => (x"4b",x"87",x"c5",x"c0"),
   346 => (x"0f",x"73",x"49",x"fd"),
   347 => (x"fa",x"c3",x"7e",x"c1"),
   348 => (x"87",x"f7",x"e1",x"49"),
   349 => (x"99",x"c2",x"49",x"70"),
   350 => (x"87",x"ea",x"c0",x"02"),
   351 => (x"bf",x"e4",x"f7",x"c2"),
   352 => (x"a8",x"b7",x"c7",x"48"),
   353 => (x"87",x"c9",x"c0",x"03"),
   354 => (x"48",x"e4",x"f7",x"c2"),
   355 => (x"d3",x"c0",x"78",x"c7"),
   356 => (x"48",x"66",x"c4",x"87"),
   357 => (x"70",x"80",x"e0",x"c1"),
   358 => (x"02",x"bf",x"6e",x"7e"),
   359 => (x"4b",x"87",x"c5",x"c0"),
   360 => (x"0f",x"73",x"49",x"fc"),
   361 => (x"48",x"75",x"7e",x"c1"),
   362 => (x"cc",x"98",x"f0",x"c3"),
   363 => (x"98",x"70",x"58",x"a6"),
   364 => (x"87",x"ce",x"c0",x"05"),
   365 => (x"e0",x"49",x"da",x"c1"),
   366 => (x"49",x"70",x"87",x"f1"),
   367 => (x"c1",x"02",x"99",x"c2"),
   368 => (x"e8",x"cf",x"87",x"f9"),
   369 => (x"87",x"d0",x"c3",x"49"),
   370 => (x"f7",x"c2",x"4b",x"70"),
   371 => (x"50",x"c0",x"48",x"dc"),
   372 => (x"97",x"dc",x"f7",x"c2"),
   373 => (x"d2",x"c1",x"05",x"bf"),
   374 => (x"05",x"66",x"c8",x"87"),
   375 => (x"c1",x"87",x"cc",x"c0"),
   376 => (x"c6",x"e0",x"49",x"da"),
   377 => (x"02",x"98",x"70",x"87"),
   378 => (x"e8",x"87",x"c0",x"c1"),
   379 => (x"c3",x"49",x"4d",x"bf"),
   380 => (x"b7",x"c8",x"99",x"ff"),
   381 => (x"ff",x"b5",x"71",x"2d"),
   382 => (x"73",x"87",x"f3",x"da"),
   383 => (x"87",x"e4",x"c2",x"49"),
   384 => (x"c0",x"02",x"98",x"70"),
   385 => (x"f7",x"c2",x"87",x"c6"),
   386 => (x"50",x"c1",x"48",x"dc"),
   387 => (x"97",x"dc",x"f7",x"c2"),
   388 => (x"d6",x"c0",x"05",x"bf"),
   389 => (x"c3",x"49",x"75",x"87"),
   390 => (x"ff",x"05",x"99",x"f0"),
   391 => (x"da",x"c1",x"87",x"cd"),
   392 => (x"c6",x"df",x"ff",x"49"),
   393 => (x"05",x"98",x"70",x"87"),
   394 => (x"c2",x"87",x"c0",x"ff"),
   395 => (x"49",x"bf",x"e4",x"f7"),
   396 => (x"c4",x"93",x"cc",x"4b"),
   397 => (x"4b",x"6b",x"83",x"66"),
   398 => (x"74",x"0f",x"73",x"71"),
   399 => (x"e9",x"c0",x"02",x"9c"),
   400 => (x"c0",x"02",x"6c",x"87"),
   401 => (x"49",x"6c",x"87",x"e4"),
   402 => (x"87",x"df",x"de",x"ff"),
   403 => (x"99",x"c1",x"49",x"70"),
   404 => (x"87",x"cb",x"c0",x"02"),
   405 => (x"c2",x"4b",x"a4",x"c4"),
   406 => (x"49",x"bf",x"e4",x"f7"),
   407 => (x"c8",x"0f",x"4b",x"6b"),
   408 => (x"c5",x"c0",x"02",x"84"),
   409 => (x"ff",x"05",x"6c",x"87"),
   410 => (x"02",x"6e",x"87",x"dc"),
   411 => (x"c2",x"87",x"c8",x"c0"),
   412 => (x"49",x"bf",x"e4",x"f7"),
   413 => (x"f4",x"87",x"e9",x"f1"),
   414 => (x"26",x"4d",x"26",x"8e"),
   415 => (x"26",x"4b",x"26",x"4c"),
   416 => (x"00",x"00",x"00",x"4f"),
   417 => (x"00",x"00",x"00",x"10"),
   418 => (x"00",x"00",x"00",x"00"),
   419 => (x"00",x"00",x"00",x"00"),
   420 => (x"00",x"00",x"00",x"00"),
   421 => (x"00",x"00",x"00",x"00"),
   422 => (x"ff",x"4a",x"71",x"1e"),
   423 => (x"72",x"49",x"bf",x"c8"),
   424 => (x"4f",x"26",x"48",x"a1"),
   425 => (x"bf",x"c8",x"ff",x"1e"),
   426 => (x"c0",x"c0",x"fe",x"89"),
   427 => (x"a9",x"c0",x"c0",x"c0"),
   428 => (x"c0",x"87",x"c4",x"01"),
   429 => (x"c1",x"87",x"c2",x"4a"),
   430 => (x"26",x"48",x"72",x"4a"),
   431 => (x"5b",x"5e",x"0e",x"4f"),
   432 => (x"71",x"0e",x"5d",x"5c"),
   433 => (x"4c",x"d4",x"ff",x"4b"),
   434 => (x"c0",x"48",x"66",x"d0"),
   435 => (x"ff",x"49",x"d6",x"78"),
   436 => (x"c3",x"87",x"d5",x"dd"),
   437 => (x"49",x"6c",x"7c",x"ff"),
   438 => (x"71",x"99",x"ff",x"c3"),
   439 => (x"f0",x"c3",x"49",x"4d"),
   440 => (x"a9",x"e0",x"c1",x"99"),
   441 => (x"c3",x"87",x"cb",x"05"),
   442 => (x"48",x"6c",x"7c",x"ff"),
   443 => (x"66",x"d0",x"98",x"c3"),
   444 => (x"ff",x"c3",x"78",x"08"),
   445 => (x"49",x"4a",x"6c",x"7c"),
   446 => (x"ff",x"c3",x"31",x"c8"),
   447 => (x"71",x"4a",x"6c",x"7c"),
   448 => (x"c8",x"49",x"72",x"b2"),
   449 => (x"7c",x"ff",x"c3",x"31"),
   450 => (x"b2",x"71",x"4a",x"6c"),
   451 => (x"31",x"c8",x"49",x"72"),
   452 => (x"6c",x"7c",x"ff",x"c3"),
   453 => (x"ff",x"b2",x"71",x"4a"),
   454 => (x"e0",x"c0",x"48",x"d0"),
   455 => (x"02",x"9b",x"73",x"78"),
   456 => (x"7b",x"72",x"87",x"c2"),
   457 => (x"4d",x"26",x"48",x"75"),
   458 => (x"4b",x"26",x"4c",x"26"),
   459 => (x"26",x"1e",x"4f",x"26"),
   460 => (x"5b",x"5e",x"0e",x"4f"),
   461 => (x"86",x"f8",x"0e",x"5c"),
   462 => (x"a6",x"c8",x"1e",x"76"),
   463 => (x"87",x"fd",x"fd",x"49"),
   464 => (x"4b",x"70",x"86",x"c4"),
   465 => (x"a8",x"c4",x"48",x"6e"),
   466 => (x"87",x"fb",x"c2",x"03"),
   467 => (x"f0",x"c3",x"4a",x"73"),
   468 => (x"aa",x"d0",x"c1",x"9a"),
   469 => (x"c1",x"87",x"c7",x"02"),
   470 => (x"c2",x"05",x"aa",x"e0"),
   471 => (x"49",x"73",x"87",x"e9"),
   472 => (x"c3",x"02",x"99",x"c8"),
   473 => (x"87",x"c6",x"ff",x"87"),
   474 => (x"9c",x"c3",x"4c",x"73"),
   475 => (x"c1",x"05",x"ac",x"c2"),
   476 => (x"66",x"c4",x"87",x"c4"),
   477 => (x"71",x"31",x"c9",x"49"),
   478 => (x"4a",x"66",x"c4",x"1e"),
   479 => (x"c2",x"92",x"cc",x"c1"),
   480 => (x"72",x"49",x"ec",x"f7"),
   481 => (x"c1",x"cd",x"fe",x"81"),
   482 => (x"ff",x"49",x"d8",x"87"),
   483 => (x"c8",x"87",x"d9",x"da"),
   484 => (x"e4",x"c2",x"1e",x"c0"),
   485 => (x"e6",x"fd",x"49",x"e4"),
   486 => (x"d0",x"ff",x"87",x"d9"),
   487 => (x"78",x"e0",x"c0",x"48"),
   488 => (x"1e",x"e4",x"e4",x"c2"),
   489 => (x"c1",x"4a",x"66",x"cc"),
   490 => (x"f7",x"c2",x"92",x"cc"),
   491 => (x"81",x"72",x"49",x"ec"),
   492 => (x"87",x"d7",x"cb",x"fe"),
   493 => (x"ac",x"c1",x"86",x"cc"),
   494 => (x"87",x"cb",x"c1",x"05"),
   495 => (x"fd",x"49",x"ee",x"c0"),
   496 => (x"c4",x"87",x"c9",x"e3"),
   497 => (x"31",x"c9",x"49",x"66"),
   498 => (x"66",x"c4",x"1e",x"71"),
   499 => (x"92",x"cc",x"c1",x"4a"),
   500 => (x"49",x"ec",x"f7",x"c2"),
   501 => (x"cb",x"fe",x"81",x"72"),
   502 => (x"e4",x"c2",x"87",x"f0"),
   503 => (x"66",x"c8",x"1e",x"e4"),
   504 => (x"92",x"cc",x"c1",x"4a"),
   505 => (x"49",x"ec",x"f7",x"c2"),
   506 => (x"c9",x"fe",x"81",x"72"),
   507 => (x"49",x"d7",x"87",x"de"),
   508 => (x"87",x"f4",x"d8",x"ff"),
   509 => (x"c2",x"1e",x"c0",x"c8"),
   510 => (x"fd",x"49",x"e4",x"e4"),
   511 => (x"cc",x"87",x"d1",x"e4"),
   512 => (x"48",x"d0",x"ff",x"86"),
   513 => (x"f8",x"78",x"e0",x"c0"),
   514 => (x"26",x"4c",x"26",x"8e"),
   515 => (x"1e",x"4f",x"26",x"4b"),
   516 => (x"b7",x"c4",x"4a",x"71"),
   517 => (x"87",x"ce",x"03",x"aa"),
   518 => (x"cc",x"c1",x"49",x"72"),
   519 => (x"ec",x"f7",x"c2",x"91"),
   520 => (x"81",x"c8",x"c1",x"81"),
   521 => (x"4f",x"26",x"79",x"c0"),
   522 => (x"5c",x"5b",x"5e",x"0e"),
   523 => (x"86",x"fc",x"0e",x"5d"),
   524 => (x"d4",x"ff",x"4a",x"71"),
   525 => (x"d4",x"4c",x"c0",x"4b"),
   526 => (x"b7",x"c3",x"4d",x"66"),
   527 => (x"c2",x"c2",x"01",x"ad"),
   528 => (x"02",x"9a",x"72",x"87"),
   529 => (x"1e",x"87",x"ec",x"c0"),
   530 => (x"cc",x"c1",x"49",x"75"),
   531 => (x"ec",x"f7",x"c2",x"91"),
   532 => (x"c8",x"80",x"71",x"48"),
   533 => (x"66",x"c4",x"58",x"a6"),
   534 => (x"fb",x"c2",x"fe",x"49"),
   535 => (x"70",x"86",x"c4",x"87"),
   536 => (x"87",x"d4",x"02",x"98"),
   537 => (x"c8",x"c1",x"49",x"6e"),
   538 => (x"6e",x"79",x"c1",x"81"),
   539 => (x"69",x"81",x"c8",x"49"),
   540 => (x"75",x"87",x"c5",x"4c"),
   541 => (x"87",x"d7",x"fe",x"49"),
   542 => (x"c8",x"48",x"d0",x"ff"),
   543 => (x"7b",x"dd",x"78",x"e1"),
   544 => (x"ff",x"c3",x"48",x"74"),
   545 => (x"74",x"7b",x"70",x"98"),
   546 => (x"29",x"b7",x"c8",x"49"),
   547 => (x"ff",x"c3",x"48",x"71"),
   548 => (x"74",x"7b",x"70",x"98"),
   549 => (x"29",x"b7",x"d0",x"49"),
   550 => (x"ff",x"c3",x"48",x"71"),
   551 => (x"74",x"7b",x"70",x"98"),
   552 => (x"28",x"b7",x"d8",x"48"),
   553 => (x"7b",x"c0",x"7b",x"70"),
   554 => (x"7b",x"7b",x"7b",x"7b"),
   555 => (x"7b",x"7b",x"7b",x"7b"),
   556 => (x"ff",x"7b",x"7b",x"7b"),
   557 => (x"e0",x"c0",x"48",x"d0"),
   558 => (x"dc",x"1e",x"75",x"78"),
   559 => (x"cc",x"d6",x"ff",x"49"),
   560 => (x"fc",x"86",x"c4",x"87"),
   561 => (x"26",x"4d",x"26",x"8e"),
   562 => (x"26",x"4b",x"26",x"4c"),
   563 => (x"00",x"00",x"00",x"4f"),
   564 => (x"ff",x"ff",x"ff",x"ff"),
   565 => (x"ff",x"ff",x"ff",x"ff"),
   566 => (x"ff",x"ff",x"ff",x"ff"),
   567 => (x"ff",x"ff",x"ff",x"ff"),
   568 => (x"00",x"00",x"28",x"e4"),
   569 => (x"33",x"49",x"56",x"53"),
   570 => (x"20",x"20",x"38",x"32"),
   571 => (x"00",x"4d",x"4f",x"52"),
   572 => (x"00",x"00",x"1b",x"d3"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

