
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"f8",x"ce",x"c3",x"87"),
    12 => (x"86",x"c0",x"c6",x"4e"),
    13 => (x"49",x"f8",x"ce",x"c3"),
    14 => (x"48",x"d0",x"fb",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"ff",x"e0"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"4a",x"66",x"c4",x"1e"),
    47 => (x"51",x"12",x"48",x"71"),
    48 => (x"26",x"87",x"fb",x"05"),
    49 => (x"48",x"73",x"1e",x"4f"),
    50 => (x"05",x"a9",x"73",x"81"),
    51 => (x"87",x"f9",x"53",x"72"),
    52 => (x"73",x"1e",x"4f",x"26"),
    53 => (x"02",x"9a",x"72",x"1e"),
    54 => (x"c0",x"87",x"e7",x"c0"),
    55 => (x"72",x"4b",x"c1",x"48"),
    56 => (x"87",x"d1",x"06",x"a9"),
    57 => (x"c9",x"06",x"82",x"72"),
    58 => (x"72",x"83",x"73",x"87"),
    59 => (x"87",x"f4",x"01",x"a9"),
    60 => (x"b2",x"c1",x"87",x"c3"),
    61 => (x"03",x"a9",x"72",x"3a"),
    62 => (x"07",x"80",x"73",x"89"),
    63 => (x"05",x"2b",x"2a",x"c1"),
    64 => (x"4b",x"26",x"87",x"f3"),
    65 => (x"75",x"1e",x"4f",x"26"),
    66 => (x"71",x"4d",x"c4",x"1e"),
    67 => (x"ff",x"04",x"a1",x"b7"),
    68 => (x"c3",x"81",x"c1",x"b9"),
    69 => (x"b7",x"72",x"07",x"bd"),
    70 => (x"ba",x"ff",x"04",x"a2"),
    71 => (x"bd",x"c1",x"82",x"c1"),
    72 => (x"87",x"ee",x"fe",x"07"),
    73 => (x"ff",x"04",x"2d",x"c1"),
    74 => (x"07",x"80",x"c1",x"b8"),
    75 => (x"b9",x"ff",x"04",x"2d"),
    76 => (x"26",x"07",x"81",x"c1"),
    77 => (x"1e",x"4f",x"26",x"4d"),
    78 => (x"c3",x"48",x"d4",x"ff"),
    79 => (x"51",x"68",x"78",x"ff"),
    80 => (x"c1",x"48",x"66",x"c4"),
    81 => (x"58",x"a6",x"c8",x"88"),
    82 => (x"eb",x"05",x"98",x"70"),
    83 => (x"1e",x"4f",x"26",x"87"),
    84 => (x"d4",x"ff",x"1e",x"73"),
    85 => (x"7b",x"ff",x"c3",x"4b"),
    86 => (x"ff",x"c3",x"4a",x"6b"),
    87 => (x"c8",x"49",x"6b",x"7b"),
    88 => (x"c3",x"b1",x"72",x"32"),
    89 => (x"4a",x"6b",x"7b",x"ff"),
    90 => (x"b2",x"71",x"31",x"c8"),
    91 => (x"6b",x"7b",x"ff",x"c3"),
    92 => (x"72",x"32",x"c8",x"49"),
    93 => (x"c4",x"48",x"71",x"b1"),
    94 => (x"26",x"4d",x"26",x"87"),
    95 => (x"26",x"4b",x"26",x"4c"),
    96 => (x"5b",x"5e",x"0e",x"4f"),
    97 => (x"71",x"0e",x"5d",x"5c"),
    98 => (x"4c",x"d4",x"ff",x"4a"),
    99 => (x"ff",x"c3",x"49",x"72"),
   100 => (x"c2",x"7c",x"71",x"99"),
   101 => (x"05",x"bf",x"d0",x"fb"),
   102 => (x"66",x"d0",x"87",x"c8"),
   103 => (x"d4",x"30",x"c9",x"48"),
   104 => (x"66",x"d0",x"58",x"a6"),
   105 => (x"c3",x"29",x"d8",x"49"),
   106 => (x"7c",x"71",x"99",x"ff"),
   107 => (x"d0",x"49",x"66",x"d0"),
   108 => (x"99",x"ff",x"c3",x"29"),
   109 => (x"66",x"d0",x"7c",x"71"),
   110 => (x"c3",x"29",x"c8",x"49"),
   111 => (x"7c",x"71",x"99",x"ff"),
   112 => (x"c3",x"49",x"66",x"d0"),
   113 => (x"7c",x"71",x"99",x"ff"),
   114 => (x"29",x"d0",x"49",x"72"),
   115 => (x"71",x"99",x"ff",x"c3"),
   116 => (x"c9",x"4b",x"6c",x"7c"),
   117 => (x"c3",x"4d",x"ff",x"f0"),
   118 => (x"d0",x"05",x"ab",x"ff"),
   119 => (x"7c",x"ff",x"c3",x"87"),
   120 => (x"8d",x"c1",x"4b",x"6c"),
   121 => (x"c3",x"87",x"c6",x"02"),
   122 => (x"f0",x"02",x"ab",x"ff"),
   123 => (x"fe",x"48",x"73",x"87"),
   124 => (x"c0",x"1e",x"87",x"c7"),
   125 => (x"48",x"d4",x"ff",x"49"),
   126 => (x"c1",x"78",x"ff",x"c3"),
   127 => (x"b7",x"c8",x"c3",x"81"),
   128 => (x"87",x"f1",x"04",x"a9"),
   129 => (x"73",x"1e",x"4f",x"26"),
   130 => (x"c4",x"87",x"e7",x"1e"),
   131 => (x"c0",x"4b",x"df",x"f8"),
   132 => (x"f0",x"ff",x"c0",x"1e"),
   133 => (x"fd",x"49",x"f7",x"c1"),
   134 => (x"86",x"c4",x"87",x"e7"),
   135 => (x"c0",x"05",x"a8",x"c1"),
   136 => (x"d4",x"ff",x"87",x"ea"),
   137 => (x"78",x"ff",x"c3",x"48"),
   138 => (x"c0",x"c0",x"c0",x"c1"),
   139 => (x"c0",x"1e",x"c0",x"c0"),
   140 => (x"e9",x"c1",x"f0",x"e1"),
   141 => (x"87",x"c9",x"fd",x"49"),
   142 => (x"98",x"70",x"86",x"c4"),
   143 => (x"ff",x"87",x"ca",x"05"),
   144 => (x"ff",x"c3",x"48",x"d4"),
   145 => (x"cb",x"48",x"c1",x"78"),
   146 => (x"87",x"e6",x"fe",x"87"),
   147 => (x"fe",x"05",x"8b",x"c1"),
   148 => (x"48",x"c0",x"87",x"fd"),
   149 => (x"1e",x"87",x"e6",x"fc"),
   150 => (x"d4",x"ff",x"1e",x"73"),
   151 => (x"78",x"ff",x"c3",x"48"),
   152 => (x"1e",x"c0",x"4b",x"d3"),
   153 => (x"c1",x"f0",x"ff",x"c0"),
   154 => (x"d4",x"fc",x"49",x"c1"),
   155 => (x"70",x"86",x"c4",x"87"),
   156 => (x"87",x"ca",x"05",x"98"),
   157 => (x"c3",x"48",x"d4",x"ff"),
   158 => (x"48",x"c1",x"78",x"ff"),
   159 => (x"f1",x"fd",x"87",x"cb"),
   160 => (x"05",x"8b",x"c1",x"87"),
   161 => (x"c0",x"87",x"db",x"ff"),
   162 => (x"87",x"f1",x"fb",x"48"),
   163 => (x"5c",x"5b",x"5e",x"0e"),
   164 => (x"4c",x"d4",x"ff",x"0e"),
   165 => (x"c6",x"87",x"db",x"fd"),
   166 => (x"e1",x"c0",x"1e",x"ea"),
   167 => (x"49",x"c8",x"c1",x"f0"),
   168 => (x"c4",x"87",x"de",x"fb"),
   169 => (x"02",x"a8",x"c1",x"86"),
   170 => (x"ea",x"fe",x"87",x"c8"),
   171 => (x"c1",x"48",x"c0",x"87"),
   172 => (x"da",x"fa",x"87",x"e2"),
   173 => (x"cf",x"49",x"70",x"87"),
   174 => (x"c6",x"99",x"ff",x"ff"),
   175 => (x"c8",x"02",x"a9",x"ea"),
   176 => (x"87",x"d3",x"fe",x"87"),
   177 => (x"cb",x"c1",x"48",x"c0"),
   178 => (x"7c",x"ff",x"c3",x"87"),
   179 => (x"fc",x"4b",x"f1",x"c0"),
   180 => (x"98",x"70",x"87",x"f4"),
   181 => (x"87",x"eb",x"c0",x"02"),
   182 => (x"ff",x"c0",x"1e",x"c0"),
   183 => (x"49",x"fa",x"c1",x"f0"),
   184 => (x"c4",x"87",x"de",x"fa"),
   185 => (x"05",x"98",x"70",x"86"),
   186 => (x"ff",x"c3",x"87",x"d9"),
   187 => (x"c3",x"49",x"6c",x"7c"),
   188 => (x"7c",x"7c",x"7c",x"ff"),
   189 => (x"99",x"c0",x"c1",x"7c"),
   190 => (x"c1",x"87",x"c4",x"02"),
   191 => (x"c0",x"87",x"d5",x"48"),
   192 => (x"c2",x"87",x"d1",x"48"),
   193 => (x"87",x"c4",x"05",x"ab"),
   194 => (x"87",x"c8",x"48",x"c0"),
   195 => (x"fe",x"05",x"8b",x"c1"),
   196 => (x"48",x"c0",x"87",x"fd"),
   197 => (x"1e",x"87",x"e4",x"f9"),
   198 => (x"fb",x"c2",x"1e",x"73"),
   199 => (x"78",x"c1",x"48",x"d0"),
   200 => (x"d0",x"ff",x"4b",x"c7"),
   201 => (x"fb",x"78",x"c2",x"48"),
   202 => (x"d0",x"ff",x"87",x"c8"),
   203 => (x"c0",x"78",x"c3",x"48"),
   204 => (x"d0",x"e5",x"c0",x"1e"),
   205 => (x"f9",x"49",x"c0",x"c1"),
   206 => (x"86",x"c4",x"87",x"c7"),
   207 => (x"c1",x"05",x"a8",x"c1"),
   208 => (x"ab",x"c2",x"4b",x"87"),
   209 => (x"c0",x"87",x"c5",x"05"),
   210 => (x"87",x"f9",x"c0",x"48"),
   211 => (x"ff",x"05",x"8b",x"c1"),
   212 => (x"f7",x"fc",x"87",x"d0"),
   213 => (x"d4",x"fb",x"c2",x"87"),
   214 => (x"05",x"98",x"70",x"58"),
   215 => (x"1e",x"c1",x"87",x"cd"),
   216 => (x"c1",x"f0",x"ff",x"c0"),
   217 => (x"d8",x"f8",x"49",x"d0"),
   218 => (x"ff",x"86",x"c4",x"87"),
   219 => (x"ff",x"c3",x"48",x"d4"),
   220 => (x"87",x"fe",x"c2",x"78"),
   221 => (x"58",x"d8",x"fb",x"c2"),
   222 => (x"c2",x"48",x"d0",x"ff"),
   223 => (x"48",x"d4",x"ff",x"78"),
   224 => (x"c1",x"78",x"ff",x"c3"),
   225 => (x"87",x"f5",x"f7",x"48"),
   226 => (x"4a",x"d4",x"ff",x"1e"),
   227 => (x"c4",x"48",x"d0",x"ff"),
   228 => (x"ff",x"c3",x"78",x"d1"),
   229 => (x"05",x"89",x"c1",x"7a"),
   230 => (x"4f",x"26",x"87",x"f8"),
   231 => (x"71",x"1e",x"73",x"1e"),
   232 => (x"cd",x"ee",x"c5",x"4b"),
   233 => (x"d4",x"ff",x"4a",x"df"),
   234 => (x"78",x"ff",x"c3",x"48"),
   235 => (x"fe",x"c3",x"48",x"68"),
   236 => (x"87",x"c5",x"02",x"a8"),
   237 => (x"ed",x"05",x"8a",x"c1"),
   238 => (x"05",x"9a",x"72",x"87"),
   239 => (x"48",x"c0",x"87",x"c5"),
   240 => (x"73",x"87",x"ea",x"c0"),
   241 => (x"87",x"cc",x"02",x"9b"),
   242 => (x"73",x"1e",x"66",x"c8"),
   243 => (x"87",x"e7",x"f5",x"49"),
   244 => (x"87",x"c6",x"86",x"c4"),
   245 => (x"fe",x"49",x"66",x"c8"),
   246 => (x"d4",x"ff",x"87",x"ee"),
   247 => (x"78",x"ff",x"c3",x"48"),
   248 => (x"05",x"9b",x"73",x"78"),
   249 => (x"d0",x"ff",x"87",x"c5"),
   250 => (x"c1",x"78",x"d0",x"48"),
   251 => (x"87",x"cd",x"f6",x"48"),
   252 => (x"71",x"1e",x"73",x"1e"),
   253 => (x"ff",x"4b",x"c0",x"4a"),
   254 => (x"ff",x"c3",x"48",x"d4"),
   255 => (x"48",x"d0",x"ff",x"78"),
   256 => (x"ff",x"78",x"c3",x"c4"),
   257 => (x"ff",x"c3",x"48",x"d4"),
   258 => (x"c0",x"1e",x"72",x"78"),
   259 => (x"d1",x"c1",x"f0",x"ff"),
   260 => (x"87",x"ed",x"f5",x"49"),
   261 => (x"98",x"70",x"86",x"c4"),
   262 => (x"c8",x"87",x"cd",x"05"),
   263 => (x"66",x"cc",x"1e",x"c0"),
   264 => (x"87",x"f8",x"fd",x"49"),
   265 => (x"4b",x"70",x"86",x"c4"),
   266 => (x"c2",x"48",x"d0",x"ff"),
   267 => (x"f5",x"48",x"73",x"78"),
   268 => (x"5e",x"0e",x"87",x"cb"),
   269 => (x"0e",x"5d",x"5c",x"5b"),
   270 => (x"ff",x"c0",x"1e",x"c0"),
   271 => (x"49",x"c9",x"c1",x"f0"),
   272 => (x"d2",x"87",x"fe",x"f4"),
   273 => (x"d8",x"fb",x"c2",x"1e"),
   274 => (x"87",x"d0",x"fd",x"49"),
   275 => (x"4c",x"c0",x"86",x"c8"),
   276 => (x"b7",x"d2",x"84",x"c1"),
   277 => (x"87",x"f8",x"04",x"ac"),
   278 => (x"97",x"d8",x"fb",x"c2"),
   279 => (x"c0",x"c3",x"49",x"bf"),
   280 => (x"a9",x"c0",x"c1",x"99"),
   281 => (x"87",x"e7",x"c0",x"05"),
   282 => (x"97",x"df",x"fb",x"c2"),
   283 => (x"31",x"d0",x"49",x"bf"),
   284 => (x"97",x"e0",x"fb",x"c2"),
   285 => (x"32",x"c8",x"4a",x"bf"),
   286 => (x"fb",x"c2",x"b1",x"72"),
   287 => (x"4a",x"bf",x"97",x"e1"),
   288 => (x"cf",x"4c",x"71",x"b1"),
   289 => (x"9c",x"ff",x"ff",x"ff"),
   290 => (x"34",x"ca",x"84",x"c1"),
   291 => (x"c2",x"87",x"e7",x"c1"),
   292 => (x"bf",x"97",x"e1",x"fb"),
   293 => (x"c6",x"31",x"c1",x"49"),
   294 => (x"e2",x"fb",x"c2",x"99"),
   295 => (x"c7",x"4a",x"bf",x"97"),
   296 => (x"b1",x"72",x"2a",x"b7"),
   297 => (x"97",x"dd",x"fb",x"c2"),
   298 => (x"cf",x"4d",x"4a",x"bf"),
   299 => (x"de",x"fb",x"c2",x"9d"),
   300 => (x"c3",x"4a",x"bf",x"97"),
   301 => (x"c2",x"32",x"ca",x"9a"),
   302 => (x"bf",x"97",x"df",x"fb"),
   303 => (x"73",x"33",x"c2",x"4b"),
   304 => (x"e0",x"fb",x"c2",x"b2"),
   305 => (x"c3",x"4b",x"bf",x"97"),
   306 => (x"b7",x"c6",x"9b",x"c0"),
   307 => (x"c2",x"b2",x"73",x"2b"),
   308 => (x"71",x"48",x"c1",x"81"),
   309 => (x"c1",x"49",x"70",x"30"),
   310 => (x"70",x"30",x"75",x"48"),
   311 => (x"c1",x"4c",x"72",x"4d"),
   312 => (x"c8",x"94",x"71",x"84"),
   313 => (x"06",x"ad",x"b7",x"c0"),
   314 => (x"34",x"c1",x"87",x"cc"),
   315 => (x"c0",x"c8",x"2d",x"b7"),
   316 => (x"ff",x"01",x"ad",x"b7"),
   317 => (x"48",x"74",x"87",x"f4"),
   318 => (x"0e",x"87",x"fe",x"f1"),
   319 => (x"5d",x"5c",x"5b",x"5e"),
   320 => (x"c3",x"86",x"f8",x"0e"),
   321 => (x"c0",x"48",x"fe",x"c3"),
   322 => (x"f6",x"fb",x"c2",x"78"),
   323 => (x"fb",x"49",x"c0",x"1e"),
   324 => (x"86",x"c4",x"87",x"de"),
   325 => (x"c5",x"05",x"98",x"70"),
   326 => (x"c9",x"48",x"c0",x"87"),
   327 => (x"4d",x"c0",x"87",x"ce"),
   328 => (x"f6",x"c0",x"7e",x"c1"),
   329 => (x"c2",x"49",x"bf",x"ef"),
   330 => (x"71",x"4a",x"ec",x"fc"),
   331 => (x"f9",x"ec",x"4b",x"c8"),
   332 => (x"05",x"98",x"70",x"87"),
   333 => (x"7e",x"c0",x"87",x"c2"),
   334 => (x"bf",x"eb",x"f6",x"c0"),
   335 => (x"c8",x"fd",x"c2",x"49"),
   336 => (x"4b",x"c8",x"71",x"4a"),
   337 => (x"70",x"87",x"e3",x"ec"),
   338 => (x"87",x"c2",x"05",x"98"),
   339 => (x"02",x"6e",x"7e",x"c0"),
   340 => (x"c3",x"87",x"fd",x"c0"),
   341 => (x"4d",x"bf",x"fc",x"c2"),
   342 => (x"9f",x"f4",x"c3",x"c3"),
   343 => (x"c5",x"48",x"7e",x"bf"),
   344 => (x"05",x"a8",x"ea",x"d6"),
   345 => (x"c2",x"c3",x"87",x"c7"),
   346 => (x"ce",x"4d",x"bf",x"fc"),
   347 => (x"ca",x"48",x"6e",x"87"),
   348 => (x"02",x"a8",x"d5",x"e9"),
   349 => (x"48",x"c0",x"87",x"c5"),
   350 => (x"c2",x"87",x"f1",x"c7"),
   351 => (x"75",x"1e",x"f6",x"fb"),
   352 => (x"87",x"ec",x"f9",x"49"),
   353 => (x"98",x"70",x"86",x"c4"),
   354 => (x"c0",x"87",x"c5",x"05"),
   355 => (x"87",x"dc",x"c7",x"48"),
   356 => (x"bf",x"eb",x"f6",x"c0"),
   357 => (x"c8",x"fd",x"c2",x"49"),
   358 => (x"4b",x"c8",x"71",x"4a"),
   359 => (x"70",x"87",x"cb",x"eb"),
   360 => (x"87",x"c8",x"05",x"98"),
   361 => (x"48",x"fe",x"c3",x"c3"),
   362 => (x"87",x"da",x"78",x"c1"),
   363 => (x"bf",x"ef",x"f6",x"c0"),
   364 => (x"ec",x"fc",x"c2",x"49"),
   365 => (x"4b",x"c8",x"71",x"4a"),
   366 => (x"70",x"87",x"ef",x"ea"),
   367 => (x"c5",x"c0",x"02",x"98"),
   368 => (x"c6",x"48",x"c0",x"87"),
   369 => (x"c3",x"c3",x"87",x"e6"),
   370 => (x"49",x"bf",x"97",x"f4"),
   371 => (x"05",x"a9",x"d5",x"c1"),
   372 => (x"c3",x"87",x"cd",x"c0"),
   373 => (x"bf",x"97",x"f5",x"c3"),
   374 => (x"a9",x"ea",x"c2",x"49"),
   375 => (x"87",x"c5",x"c0",x"02"),
   376 => (x"c7",x"c6",x"48",x"c0"),
   377 => (x"f6",x"fb",x"c2",x"87"),
   378 => (x"48",x"7e",x"bf",x"97"),
   379 => (x"02",x"a8",x"e9",x"c3"),
   380 => (x"6e",x"87",x"ce",x"c0"),
   381 => (x"a8",x"eb",x"c3",x"48"),
   382 => (x"87",x"c5",x"c0",x"02"),
   383 => (x"eb",x"c5",x"48",x"c0"),
   384 => (x"c1",x"fc",x"c2",x"87"),
   385 => (x"99",x"49",x"bf",x"97"),
   386 => (x"87",x"cc",x"c0",x"05"),
   387 => (x"97",x"c2",x"fc",x"c2"),
   388 => (x"a9",x"c2",x"49",x"bf"),
   389 => (x"87",x"c5",x"c0",x"02"),
   390 => (x"cf",x"c5",x"48",x"c0"),
   391 => (x"c3",x"fc",x"c2",x"87"),
   392 => (x"c3",x"48",x"bf",x"97"),
   393 => (x"70",x"58",x"fa",x"c3"),
   394 => (x"88",x"c1",x"48",x"4c"),
   395 => (x"58",x"fe",x"c3",x"c3"),
   396 => (x"97",x"c4",x"fc",x"c2"),
   397 => (x"81",x"75",x"49",x"bf"),
   398 => (x"97",x"c5",x"fc",x"c2"),
   399 => (x"32",x"c8",x"4a",x"bf"),
   400 => (x"c3",x"7e",x"a1",x"72"),
   401 => (x"6e",x"48",x"cb",x"c8"),
   402 => (x"c6",x"fc",x"c2",x"78"),
   403 => (x"c8",x"48",x"bf",x"97"),
   404 => (x"c3",x"c3",x"58",x"a6"),
   405 => (x"c2",x"02",x"bf",x"fe"),
   406 => (x"f6",x"c0",x"87",x"d4"),
   407 => (x"c2",x"49",x"bf",x"eb"),
   408 => (x"71",x"4a",x"c8",x"fd"),
   409 => (x"c1",x"e8",x"4b",x"c8"),
   410 => (x"02",x"98",x"70",x"87"),
   411 => (x"c0",x"87",x"c5",x"c0"),
   412 => (x"87",x"f8",x"c3",x"48"),
   413 => (x"bf",x"f6",x"c3",x"c3"),
   414 => (x"df",x"c8",x"c3",x"4c"),
   415 => (x"db",x"fc",x"c2",x"5c"),
   416 => (x"c8",x"49",x"bf",x"97"),
   417 => (x"da",x"fc",x"c2",x"31"),
   418 => (x"a1",x"4a",x"bf",x"97"),
   419 => (x"dc",x"fc",x"c2",x"49"),
   420 => (x"d0",x"4a",x"bf",x"97"),
   421 => (x"49",x"a1",x"72",x"32"),
   422 => (x"97",x"dd",x"fc",x"c2"),
   423 => (x"32",x"d8",x"4a",x"bf"),
   424 => (x"c4",x"49",x"a1",x"72"),
   425 => (x"c8",x"c3",x"91",x"66"),
   426 => (x"c3",x"81",x"bf",x"cb"),
   427 => (x"c2",x"59",x"d3",x"c8"),
   428 => (x"bf",x"97",x"e3",x"fc"),
   429 => (x"c2",x"32",x"c8",x"4a"),
   430 => (x"bf",x"97",x"e2",x"fc"),
   431 => (x"c2",x"4a",x"a2",x"4b"),
   432 => (x"bf",x"97",x"e4",x"fc"),
   433 => (x"73",x"33",x"d0",x"4b"),
   434 => (x"fc",x"c2",x"4a",x"a2"),
   435 => (x"4b",x"bf",x"97",x"e5"),
   436 => (x"33",x"d8",x"9b",x"cf"),
   437 => (x"c3",x"4a",x"a2",x"73"),
   438 => (x"c3",x"5a",x"d7",x"c8"),
   439 => (x"4a",x"bf",x"d3",x"c8"),
   440 => (x"92",x"74",x"8a",x"c2"),
   441 => (x"48",x"d7",x"c8",x"c3"),
   442 => (x"c1",x"78",x"a1",x"72"),
   443 => (x"fc",x"c2",x"87",x"ca"),
   444 => (x"49",x"bf",x"97",x"c8"),
   445 => (x"fc",x"c2",x"31",x"c8"),
   446 => (x"4a",x"bf",x"97",x"c7"),
   447 => (x"c4",x"c3",x"49",x"a1"),
   448 => (x"c4",x"c3",x"59",x"c6"),
   449 => (x"c5",x"49",x"bf",x"c2"),
   450 => (x"81",x"ff",x"c7",x"31"),
   451 => (x"c8",x"c3",x"29",x"c9"),
   452 => (x"fc",x"c2",x"59",x"df"),
   453 => (x"4a",x"bf",x"97",x"cd"),
   454 => (x"fc",x"c2",x"32",x"c8"),
   455 => (x"4b",x"bf",x"97",x"cc"),
   456 => (x"66",x"c4",x"4a",x"a2"),
   457 => (x"c3",x"82",x"6e",x"92"),
   458 => (x"c3",x"5a",x"db",x"c8"),
   459 => (x"c0",x"48",x"d3",x"c8"),
   460 => (x"cf",x"c8",x"c3",x"78"),
   461 => (x"78",x"a1",x"72",x"48"),
   462 => (x"48",x"df",x"c8",x"c3"),
   463 => (x"bf",x"d3",x"c8",x"c3"),
   464 => (x"e3",x"c8",x"c3",x"78"),
   465 => (x"d7",x"c8",x"c3",x"48"),
   466 => (x"c3",x"c3",x"78",x"bf"),
   467 => (x"c0",x"02",x"bf",x"fe"),
   468 => (x"48",x"74",x"87",x"c9"),
   469 => (x"7e",x"70",x"30",x"c4"),
   470 => (x"c3",x"87",x"c9",x"c0"),
   471 => (x"48",x"bf",x"db",x"c8"),
   472 => (x"7e",x"70",x"30",x"c4"),
   473 => (x"48",x"c2",x"c4",x"c3"),
   474 => (x"48",x"c1",x"78",x"6e"),
   475 => (x"4d",x"26",x"8e",x"f8"),
   476 => (x"4b",x"26",x"4c",x"26"),
   477 => (x"5e",x"0e",x"4f",x"26"),
   478 => (x"0e",x"5d",x"5c",x"5b"),
   479 => (x"c3",x"c3",x"4a",x"71"),
   480 => (x"cb",x"02",x"bf",x"fe"),
   481 => (x"c7",x"4b",x"72",x"87"),
   482 => (x"c1",x"4c",x"72",x"2b"),
   483 => (x"87",x"c9",x"9c",x"ff"),
   484 => (x"2b",x"c8",x"4b",x"72"),
   485 => (x"ff",x"c3",x"4c",x"72"),
   486 => (x"cb",x"c8",x"c3",x"9c"),
   487 => (x"f6",x"c0",x"83",x"bf"),
   488 => (x"02",x"ab",x"bf",x"e7"),
   489 => (x"f6",x"c0",x"87",x"d9"),
   490 => (x"fb",x"c2",x"5b",x"eb"),
   491 => (x"49",x"73",x"1e",x"f6"),
   492 => (x"c4",x"87",x"fd",x"f0"),
   493 => (x"05",x"98",x"70",x"86"),
   494 => (x"48",x"c0",x"87",x"c5"),
   495 => (x"c3",x"87",x"e6",x"c0"),
   496 => (x"02",x"bf",x"fe",x"c3"),
   497 => (x"49",x"74",x"87",x"d2"),
   498 => (x"fb",x"c2",x"91",x"c4"),
   499 => (x"4d",x"69",x"81",x"f6"),
   500 => (x"ff",x"ff",x"ff",x"cf"),
   501 => (x"87",x"cb",x"9d",x"ff"),
   502 => (x"91",x"c2",x"49",x"74"),
   503 => (x"81",x"f6",x"fb",x"c2"),
   504 => (x"75",x"4d",x"69",x"9f"),
   505 => (x"87",x"c6",x"fe",x"48"),
   506 => (x"5c",x"5b",x"5e",x"0e"),
   507 => (x"71",x"1e",x"0e",x"5d"),
   508 => (x"c1",x"1e",x"c0",x"4d"),
   509 => (x"87",x"d7",x"cf",x"49"),
   510 => (x"4c",x"70",x"86",x"c4"),
   511 => (x"c0",x"c1",x"02",x"9c"),
   512 => (x"c6",x"c4",x"c3",x"87"),
   513 => (x"e1",x"49",x"75",x"4a"),
   514 => (x"98",x"70",x"87",x"c5"),
   515 => (x"87",x"f1",x"c0",x"02"),
   516 => (x"49",x"75",x"4a",x"74"),
   517 => (x"eb",x"e1",x"4b",x"cb"),
   518 => (x"02",x"98",x"70",x"87"),
   519 => (x"c0",x"87",x"e2",x"c0"),
   520 => (x"02",x"9c",x"74",x"1e"),
   521 => (x"a6",x"c4",x"87",x"c7"),
   522 => (x"c5",x"78",x"c0",x"48"),
   523 => (x"48",x"a6",x"c4",x"87"),
   524 => (x"66",x"c4",x"78",x"c1"),
   525 => (x"87",x"d7",x"ce",x"49"),
   526 => (x"4c",x"70",x"86",x"c4"),
   527 => (x"c0",x"ff",x"05",x"9c"),
   528 => (x"26",x"48",x"74",x"87"),
   529 => (x"0e",x"87",x"e7",x"fc"),
   530 => (x"5d",x"5c",x"5b",x"5e"),
   531 => (x"4b",x"71",x"1e",x"0e"),
   532 => (x"87",x"c5",x"05",x"9b"),
   533 => (x"e5",x"c1",x"48",x"c0"),
   534 => (x"4d",x"a3",x"c8",x"87"),
   535 => (x"66",x"d4",x"7d",x"c0"),
   536 => (x"d4",x"87",x"c7",x"02"),
   537 => (x"05",x"bf",x"97",x"66"),
   538 => (x"48",x"c0",x"87",x"c5"),
   539 => (x"d4",x"87",x"cf",x"c1"),
   540 => (x"f3",x"fd",x"49",x"66"),
   541 => (x"9c",x"4c",x"70",x"87"),
   542 => (x"87",x"c0",x"c1",x"02"),
   543 => (x"69",x"49",x"a4",x"dc"),
   544 => (x"49",x"a4",x"da",x"7d"),
   545 => (x"9f",x"4a",x"a3",x"c4"),
   546 => (x"c3",x"c3",x"7a",x"69"),
   547 => (x"d2",x"02",x"bf",x"fe"),
   548 => (x"49",x"a4",x"d4",x"87"),
   549 => (x"c0",x"49",x"69",x"9f"),
   550 => (x"71",x"99",x"ff",x"ff"),
   551 => (x"70",x"30",x"d0",x"48"),
   552 => (x"c0",x"87",x"c2",x"7e"),
   553 => (x"48",x"49",x"6e",x"7e"),
   554 => (x"7a",x"70",x"80",x"6a"),
   555 => (x"a3",x"cc",x"7b",x"c0"),
   556 => (x"d0",x"79",x"6a",x"49"),
   557 => (x"79",x"c0",x"49",x"a3"),
   558 => (x"87",x"c2",x"48",x"74"),
   559 => (x"fa",x"26",x"48",x"c0"),
   560 => (x"5e",x"0e",x"87",x"ec"),
   561 => (x"0e",x"5d",x"5c",x"5b"),
   562 => (x"f6",x"c0",x"4c",x"71"),
   563 => (x"78",x"ff",x"48",x"e7"),
   564 => (x"c1",x"02",x"9c",x"74"),
   565 => (x"a4",x"c8",x"87",x"ca"),
   566 => (x"c1",x"02",x"69",x"49"),
   567 => (x"66",x"d0",x"87",x"c2"),
   568 => (x"82",x"49",x"6c",x"4a"),
   569 => (x"d0",x"5a",x"a6",x"d4"),
   570 => (x"c3",x"b9",x"4d",x"66"),
   571 => (x"4a",x"bf",x"fa",x"c3"),
   572 => (x"99",x"72",x"ba",x"ff"),
   573 => (x"c0",x"02",x"99",x"71"),
   574 => (x"a4",x"c4",x"87",x"e4"),
   575 => (x"f9",x"49",x"6b",x"4b"),
   576 => (x"7b",x"70",x"87",x"f4"),
   577 => (x"bf",x"f6",x"c3",x"c3"),
   578 => (x"71",x"81",x"6c",x"49"),
   579 => (x"c3",x"b9",x"75",x"7c"),
   580 => (x"4a",x"bf",x"fa",x"c3"),
   581 => (x"99",x"72",x"ba",x"ff"),
   582 => (x"ff",x"05",x"99",x"71"),
   583 => (x"7c",x"75",x"87",x"dc"),
   584 => (x"1e",x"87",x"cb",x"f9"),
   585 => (x"4b",x"71",x"1e",x"73"),
   586 => (x"87",x"c7",x"02",x"9b"),
   587 => (x"69",x"49",x"a3",x"c8"),
   588 => (x"c0",x"87",x"c5",x"05"),
   589 => (x"87",x"eb",x"c0",x"48"),
   590 => (x"bf",x"cf",x"c8",x"c3"),
   591 => (x"49",x"a3",x"c4",x"4a"),
   592 => (x"89",x"c2",x"49",x"69"),
   593 => (x"bf",x"f6",x"c3",x"c3"),
   594 => (x"4a",x"a2",x"71",x"91"),
   595 => (x"bf",x"fa",x"c3",x"c3"),
   596 => (x"71",x"99",x"6b",x"49"),
   597 => (x"66",x"c8",x"4a",x"a2"),
   598 => (x"ea",x"49",x"72",x"1e"),
   599 => (x"86",x"c4",x"87",x"d2"),
   600 => (x"f8",x"48",x"49",x"70"),
   601 => (x"5e",x"0e",x"87",x"cc"),
   602 => (x"0e",x"5d",x"5c",x"5b"),
   603 => (x"d4",x"4b",x"71",x"1e"),
   604 => (x"2c",x"c9",x"4c",x"66"),
   605 => (x"c1",x"02",x"9b",x"73"),
   606 => (x"a3",x"c8",x"87",x"cf"),
   607 => (x"c1",x"02",x"69",x"49"),
   608 => (x"a3",x"d0",x"87",x"c7"),
   609 => (x"7d",x"66",x"d4",x"4d"),
   610 => (x"bf",x"fa",x"c3",x"c3"),
   611 => (x"6b",x"b9",x"ff",x"49"),
   612 => (x"71",x"7e",x"99",x"4a"),
   613 => (x"87",x"cd",x"03",x"ac"),
   614 => (x"cc",x"7d",x"7b",x"c0"),
   615 => (x"a3",x"c4",x"4a",x"a3"),
   616 => (x"c2",x"79",x"6a",x"49"),
   617 => (x"74",x"8c",x"72",x"87"),
   618 => (x"87",x"dd",x"02",x"9c"),
   619 => (x"49",x"73",x"1e",x"49"),
   620 => (x"c4",x"87",x"cf",x"fc"),
   621 => (x"49",x"66",x"d4",x"86"),
   622 => (x"02",x"99",x"ff",x"c7"),
   623 => (x"fb",x"c2",x"87",x"cb"),
   624 => (x"49",x"73",x"1e",x"f6"),
   625 => (x"c4",x"87",x"dc",x"fd"),
   626 => (x"e1",x"f6",x"26",x"86"),
   627 => (x"5b",x"5e",x"0e",x"87"),
   628 => (x"f0",x"0e",x"5d",x"5c"),
   629 => (x"59",x"a6",x"d0",x"86"),
   630 => (x"4b",x"66",x"e4",x"c0"),
   631 => (x"ca",x"02",x"66",x"cc"),
   632 => (x"80",x"c8",x"48",x"87"),
   633 => (x"bf",x"6e",x"7e",x"70"),
   634 => (x"c0",x"87",x"c5",x"05"),
   635 => (x"87",x"ec",x"c3",x"48"),
   636 => (x"d0",x"4c",x"66",x"cc"),
   637 => (x"c4",x"49",x"73",x"84"),
   638 => (x"78",x"6c",x"48",x"a6"),
   639 => (x"c4",x"81",x"66",x"c4"),
   640 => (x"78",x"bf",x"6e",x"80"),
   641 => (x"06",x"a9",x"66",x"c8"),
   642 => (x"c4",x"49",x"87",x"c6"),
   643 => (x"4b",x"71",x"89",x"66"),
   644 => (x"01",x"ab",x"b7",x"c0"),
   645 => (x"c3",x"48",x"87",x"c4"),
   646 => (x"66",x"c4",x"87",x"c2"),
   647 => (x"98",x"ff",x"c7",x"48"),
   648 => (x"02",x"6e",x"7e",x"70"),
   649 => (x"c8",x"87",x"c9",x"c1"),
   650 => (x"89",x"6e",x"49",x"c0"),
   651 => (x"fb",x"c2",x"4a",x"71"),
   652 => (x"85",x"6e",x"4d",x"f6"),
   653 => (x"06",x"aa",x"b7",x"73"),
   654 => (x"72",x"4a",x"87",x"c1"),
   655 => (x"66",x"c4",x"48",x"49"),
   656 => (x"72",x"7c",x"70",x"80"),
   657 => (x"8a",x"c1",x"49",x"8b"),
   658 => (x"d9",x"02",x"99",x"71"),
   659 => (x"66",x"e0",x"c0",x"87"),
   660 => (x"c0",x"50",x"15",x"48"),
   661 => (x"c1",x"48",x"66",x"e0"),
   662 => (x"a6",x"e4",x"c0",x"80"),
   663 => (x"c1",x"49",x"72",x"58"),
   664 => (x"05",x"99",x"71",x"8a"),
   665 => (x"1e",x"c1",x"87",x"e7"),
   666 => (x"f9",x"49",x"66",x"d0"),
   667 => (x"86",x"c4",x"87",x"d4"),
   668 => (x"06",x"ab",x"b7",x"c0"),
   669 => (x"c0",x"87",x"e3",x"c1"),
   670 => (x"c7",x"4d",x"66",x"e0"),
   671 => (x"06",x"ab",x"b7",x"ff"),
   672 => (x"75",x"87",x"e2",x"c0"),
   673 => (x"49",x"66",x"d0",x"1e"),
   674 => (x"c8",x"87",x"d8",x"fa"),
   675 => (x"48",x"6c",x"85",x"c0"),
   676 => (x"70",x"80",x"c0",x"c8"),
   677 => (x"8b",x"c0",x"c8",x"7c"),
   678 => (x"66",x"d4",x"1e",x"c1"),
   679 => (x"87",x"e2",x"f8",x"49"),
   680 => (x"ee",x"c0",x"86",x"c8"),
   681 => (x"f6",x"fb",x"c2",x"87"),
   682 => (x"49",x"66",x"d0",x"1e"),
   683 => (x"c4",x"87",x"f4",x"f9"),
   684 => (x"f6",x"fb",x"c2",x"86"),
   685 => (x"48",x"49",x"73",x"4a"),
   686 => (x"7c",x"70",x"80",x"6c"),
   687 => (x"8b",x"c1",x"49",x"73"),
   688 => (x"ce",x"02",x"99",x"71"),
   689 => (x"7d",x"97",x"12",x"87"),
   690 => (x"49",x"73",x"85",x"c1"),
   691 => (x"99",x"71",x"8b",x"c1"),
   692 => (x"c0",x"87",x"f2",x"05"),
   693 => (x"fe",x"01",x"ab",x"b7"),
   694 => (x"48",x"c1",x"87",x"e1"),
   695 => (x"cd",x"f2",x"8e",x"f0"),
   696 => (x"5b",x"5e",x"0e",x"87"),
   697 => (x"71",x"0e",x"5d",x"5c"),
   698 => (x"c7",x"02",x"9b",x"4b"),
   699 => (x"4d",x"a3",x"c8",x"87"),
   700 => (x"87",x"c5",x"05",x"6d"),
   701 => (x"fd",x"c0",x"48",x"ff"),
   702 => (x"4c",x"a3",x"d0",x"87"),
   703 => (x"ff",x"c7",x"49",x"6c"),
   704 => (x"87",x"d8",x"05",x"99"),
   705 => (x"87",x"c9",x"02",x"6c"),
   706 => (x"49",x"73",x"1e",x"c1"),
   707 => (x"c4",x"87",x"f3",x"f6"),
   708 => (x"f6",x"fb",x"c2",x"86"),
   709 => (x"f8",x"49",x"73",x"1e"),
   710 => (x"86",x"c4",x"87",x"c9"),
   711 => (x"aa",x"6d",x"4a",x"6c"),
   712 => (x"ff",x"87",x"c4",x"04"),
   713 => (x"c1",x"87",x"cf",x"48"),
   714 => (x"49",x"72",x"7c",x"a2"),
   715 => (x"c2",x"99",x"ff",x"c7"),
   716 => (x"97",x"81",x"f6",x"fb"),
   717 => (x"f5",x"f0",x"48",x"69"),
   718 => (x"1e",x"73",x"1e",x"87"),
   719 => (x"02",x"9b",x"4b",x"71"),
   720 => (x"c3",x"87",x"e4",x"c0"),
   721 => (x"73",x"5b",x"e3",x"c8"),
   722 => (x"c3",x"8a",x"c2",x"4a"),
   723 => (x"49",x"bf",x"f6",x"c3"),
   724 => (x"cf",x"c8",x"c3",x"92"),
   725 => (x"80",x"72",x"48",x"bf"),
   726 => (x"58",x"e7",x"c8",x"c3"),
   727 => (x"30",x"c4",x"48",x"71"),
   728 => (x"58",x"c6",x"c4",x"c3"),
   729 => (x"c3",x"87",x"ed",x"c0"),
   730 => (x"c3",x"48",x"df",x"c8"),
   731 => (x"78",x"bf",x"d3",x"c8"),
   732 => (x"48",x"e3",x"c8",x"c3"),
   733 => (x"bf",x"d7",x"c8",x"c3"),
   734 => (x"fe",x"c3",x"c3",x"78"),
   735 => (x"87",x"c9",x"02",x"bf"),
   736 => (x"bf",x"f6",x"c3",x"c3"),
   737 => (x"c7",x"31",x"c4",x"49"),
   738 => (x"db",x"c8",x"c3",x"87"),
   739 => (x"31",x"c4",x"49",x"bf"),
   740 => (x"59",x"c6",x"c4",x"c3"),
   741 => (x"0e",x"87",x"db",x"ef"),
   742 => (x"0e",x"5c",x"5b",x"5e"),
   743 => (x"4b",x"c0",x"4a",x"71"),
   744 => (x"c0",x"02",x"9a",x"72"),
   745 => (x"a2",x"da",x"87",x"e1"),
   746 => (x"4b",x"69",x"9f",x"49"),
   747 => (x"bf",x"fe",x"c3",x"c3"),
   748 => (x"d4",x"87",x"cf",x"02"),
   749 => (x"69",x"9f",x"49",x"a2"),
   750 => (x"ff",x"c0",x"4c",x"49"),
   751 => (x"34",x"d0",x"9c",x"ff"),
   752 => (x"4c",x"c0",x"87",x"c2"),
   753 => (x"73",x"b3",x"49",x"74"),
   754 => (x"87",x"ed",x"fd",x"49"),
   755 => (x"0e",x"87",x"e1",x"ee"),
   756 => (x"5d",x"5c",x"5b",x"5e"),
   757 => (x"71",x"86",x"f4",x"0e"),
   758 => (x"72",x"7e",x"c0",x"4a"),
   759 => (x"87",x"d8",x"02",x"9a"),
   760 => (x"48",x"f2",x"fb",x"c2"),
   761 => (x"fb",x"c2",x"78",x"c0"),
   762 => (x"c8",x"c3",x"48",x"ea"),
   763 => (x"c2",x"78",x"bf",x"e3"),
   764 => (x"c3",x"48",x"ee",x"fb"),
   765 => (x"78",x"bf",x"df",x"c8"),
   766 => (x"48",x"d3",x"c4",x"c3"),
   767 => (x"c4",x"c3",x"50",x"c0"),
   768 => (x"c2",x"49",x"bf",x"c2"),
   769 => (x"4a",x"bf",x"f2",x"fb"),
   770 => (x"c4",x"03",x"aa",x"71"),
   771 => (x"49",x"72",x"87",x"c0"),
   772 => (x"c0",x"05",x"99",x"cf"),
   773 => (x"fb",x"c2",x"87",x"e1"),
   774 => (x"fb",x"c2",x"1e",x"f6"),
   775 => (x"c2",x"49",x"bf",x"ea"),
   776 => (x"c1",x"48",x"ea",x"fb"),
   777 => (x"ff",x"71",x"78",x"a1"),
   778 => (x"c4",x"87",x"c5",x"df"),
   779 => (x"e3",x"f6",x"c0",x"86"),
   780 => (x"f6",x"fb",x"c2",x"48"),
   781 => (x"c0",x"87",x"cc",x"78"),
   782 => (x"48",x"bf",x"e3",x"f6"),
   783 => (x"c0",x"80",x"e0",x"c0"),
   784 => (x"c2",x"58",x"e7",x"f6"),
   785 => (x"48",x"bf",x"f2",x"fb"),
   786 => (x"fb",x"c2",x"80",x"c1"),
   787 => (x"a3",x"27",x"58",x"f6"),
   788 => (x"bf",x"00",x"00",x"0d"),
   789 => (x"9d",x"4d",x"bf",x"97"),
   790 => (x"87",x"e2",x"c2",x"02"),
   791 => (x"02",x"ad",x"e5",x"c3"),
   792 => (x"c0",x"87",x"db",x"c2"),
   793 => (x"4b",x"bf",x"e3",x"f6"),
   794 => (x"11",x"49",x"a3",x"cb"),
   795 => (x"05",x"ac",x"cf",x"4c"),
   796 => (x"75",x"87",x"d2",x"c1"),
   797 => (x"c1",x"99",x"df",x"49"),
   798 => (x"c3",x"91",x"cd",x"89"),
   799 => (x"c1",x"81",x"c6",x"c4"),
   800 => (x"51",x"12",x"4a",x"a3"),
   801 => (x"12",x"4a",x"a3",x"c3"),
   802 => (x"4a",x"a3",x"c5",x"51"),
   803 => (x"a3",x"c7",x"51",x"12"),
   804 => (x"c9",x"51",x"12",x"4a"),
   805 => (x"51",x"12",x"4a",x"a3"),
   806 => (x"12",x"4a",x"a3",x"ce"),
   807 => (x"4a",x"a3",x"d0",x"51"),
   808 => (x"a3",x"d2",x"51",x"12"),
   809 => (x"d4",x"51",x"12",x"4a"),
   810 => (x"51",x"12",x"4a",x"a3"),
   811 => (x"12",x"4a",x"a3",x"d6"),
   812 => (x"4a",x"a3",x"d8",x"51"),
   813 => (x"a3",x"dc",x"51",x"12"),
   814 => (x"de",x"51",x"12",x"4a"),
   815 => (x"51",x"12",x"4a",x"a3"),
   816 => (x"f9",x"c0",x"7e",x"c1"),
   817 => (x"c8",x"49",x"74",x"87"),
   818 => (x"ea",x"c0",x"05",x"99"),
   819 => (x"d0",x"49",x"74",x"87"),
   820 => (x"87",x"d0",x"05",x"99"),
   821 => (x"c0",x"02",x"66",x"dc"),
   822 => (x"49",x"73",x"87",x"ca"),
   823 => (x"70",x"0f",x"66",x"dc"),
   824 => (x"87",x"d3",x"02",x"98"),
   825 => (x"c6",x"c0",x"05",x"6e"),
   826 => (x"c6",x"c4",x"c3",x"87"),
   827 => (x"c0",x"50",x"c0",x"48"),
   828 => (x"48",x"bf",x"e3",x"f6"),
   829 => (x"c3",x"87",x"e7",x"c2"),
   830 => (x"c0",x"48",x"d3",x"c4"),
   831 => (x"c4",x"c3",x"7e",x"50"),
   832 => (x"c2",x"49",x"bf",x"c2"),
   833 => (x"4a",x"bf",x"f2",x"fb"),
   834 => (x"fc",x"04",x"aa",x"71"),
   835 => (x"c8",x"c3",x"87",x"c0"),
   836 => (x"c0",x"05",x"bf",x"e3"),
   837 => (x"c3",x"c3",x"87",x"c8"),
   838 => (x"c1",x"02",x"bf",x"fe"),
   839 => (x"f6",x"c0",x"87",x"fe"),
   840 => (x"78",x"ff",x"48",x"e7"),
   841 => (x"bf",x"ee",x"fb",x"c2"),
   842 => (x"87",x"ca",x"e9",x"49"),
   843 => (x"fb",x"c2",x"49",x"70"),
   844 => (x"a6",x"c4",x"59",x"f2"),
   845 => (x"ee",x"fb",x"c2",x"48"),
   846 => (x"c3",x"c3",x"78",x"bf"),
   847 => (x"c0",x"02",x"bf",x"fe"),
   848 => (x"66",x"c4",x"87",x"d8"),
   849 => (x"ff",x"ff",x"cf",x"49"),
   850 => (x"a9",x"99",x"f8",x"ff"),
   851 => (x"87",x"c5",x"c0",x"02"),
   852 => (x"e1",x"c0",x"4d",x"c0"),
   853 => (x"c0",x"4d",x"c1",x"87"),
   854 => (x"66",x"c4",x"87",x"dc"),
   855 => (x"f8",x"ff",x"cf",x"49"),
   856 => (x"c0",x"02",x"a9",x"99"),
   857 => (x"a6",x"c8",x"87",x"c8"),
   858 => (x"c0",x"78",x"c0",x"48"),
   859 => (x"a6",x"c8",x"87",x"c5"),
   860 => (x"c8",x"78",x"c1",x"48"),
   861 => (x"9d",x"75",x"4d",x"66"),
   862 => (x"87",x"e0",x"c0",x"05"),
   863 => (x"c2",x"49",x"66",x"c4"),
   864 => (x"f6",x"c3",x"c3",x"89"),
   865 => (x"c3",x"91",x"4a",x"bf"),
   866 => (x"4a",x"bf",x"cf",x"c8"),
   867 => (x"48",x"ea",x"fb",x"c2"),
   868 => (x"c2",x"78",x"a1",x"72"),
   869 => (x"c0",x"48",x"f2",x"fb"),
   870 => (x"87",x"e2",x"f9",x"78"),
   871 => (x"8e",x"f4",x"48",x"c0"),
   872 => (x"00",x"87",x"cb",x"e7"),
   873 => (x"ff",x"00",x"00",x"00"),
   874 => (x"b3",x"ff",x"ff",x"ff"),
   875 => (x"bc",x"00",x"00",x"0d"),
   876 => (x"46",x"00",x"00",x"0d"),
   877 => (x"32",x"33",x"54",x"41"),
   878 => (x"00",x"20",x"20",x"20"),
   879 => (x"31",x"54",x"41",x"46"),
   880 => (x"20",x"20",x"20",x"36"),
   881 => (x"c8",x"c3",x"1e",x"00"),
   882 => (x"dd",x"48",x"bf",x"e8"),
   883 => (x"87",x"c9",x"05",x"a8"),
   884 => (x"87",x"e8",x"fd",x"c0"),
   885 => (x"c8",x"4a",x"49",x"70"),
   886 => (x"48",x"d4",x"ff",x"87"),
   887 => (x"68",x"78",x"ff",x"c3"),
   888 => (x"26",x"48",x"72",x"4a"),
   889 => (x"c8",x"c3",x"1e",x"4f"),
   890 => (x"dd",x"48",x"bf",x"e8"),
   891 => (x"87",x"c6",x"05",x"a8"),
   892 => (x"87",x"f4",x"fc",x"c0"),
   893 => (x"d4",x"ff",x"87",x"d9"),
   894 => (x"78",x"ff",x"c3",x"48"),
   895 => (x"c8",x"48",x"d0",x"ff"),
   896 => (x"d4",x"ff",x"78",x"e1"),
   897 => (x"c3",x"78",x"d4",x"48"),
   898 => (x"ff",x"48",x"e7",x"c8"),
   899 => (x"26",x"50",x"bf",x"d4"),
   900 => (x"d0",x"ff",x"1e",x"4f"),
   901 => (x"78",x"e0",x"c0",x"48"),
   902 => (x"fe",x"1e",x"4f",x"26"),
   903 => (x"49",x"70",x"87",x"e7"),
   904 => (x"87",x"c6",x"02",x"99"),
   905 => (x"05",x"a9",x"fb",x"c0"),
   906 => (x"48",x"71",x"87",x"f1"),
   907 => (x"5e",x"0e",x"4f",x"26"),
   908 => (x"71",x"0e",x"5c",x"5b"),
   909 => (x"fe",x"4c",x"c0",x"4b"),
   910 => (x"49",x"70",x"87",x"cb"),
   911 => (x"f9",x"c0",x"02",x"99"),
   912 => (x"a9",x"ec",x"c0",x"87"),
   913 => (x"87",x"f2",x"c0",x"02"),
   914 => (x"02",x"a9",x"fb",x"c0"),
   915 => (x"cc",x"87",x"eb",x"c0"),
   916 => (x"03",x"ac",x"b7",x"66"),
   917 => (x"66",x"d0",x"87",x"c7"),
   918 => (x"71",x"87",x"c2",x"02"),
   919 => (x"02",x"99",x"71",x"53"),
   920 => (x"84",x"c1",x"87",x"c2"),
   921 => (x"70",x"87",x"de",x"fd"),
   922 => (x"cd",x"02",x"99",x"49"),
   923 => (x"a9",x"ec",x"c0",x"87"),
   924 => (x"c0",x"87",x"c7",x"02"),
   925 => (x"ff",x"05",x"a9",x"fb"),
   926 => (x"66",x"d0",x"87",x"d5"),
   927 => (x"c0",x"87",x"c3",x"02"),
   928 => (x"ec",x"c0",x"7b",x"97"),
   929 => (x"87",x"c4",x"05",x"a9"),
   930 => (x"87",x"c5",x"4a",x"74"),
   931 => (x"0a",x"c0",x"4a",x"74"),
   932 => (x"c2",x"48",x"72",x"8a"),
   933 => (x"26",x"4d",x"26",x"87"),
   934 => (x"26",x"4b",x"26",x"4c"),
   935 => (x"e4",x"fc",x"1e",x"4f"),
   936 => (x"c0",x"49",x"70",x"87"),
   937 => (x"04",x"a9",x"b7",x"f0"),
   938 => (x"f9",x"c0",x"87",x"ca"),
   939 => (x"c3",x"01",x"a9",x"b7"),
   940 => (x"89",x"f0",x"c0",x"87"),
   941 => (x"a9",x"b7",x"c1",x"c1"),
   942 => (x"c1",x"87",x"ca",x"04"),
   943 => (x"01",x"a9",x"b7",x"da"),
   944 => (x"f7",x"c0",x"87",x"c3"),
   945 => (x"26",x"48",x"71",x"89"),
   946 => (x"5b",x"5e",x"0e",x"4f"),
   947 => (x"4a",x"71",x"0e",x"5c"),
   948 => (x"72",x"4c",x"d4",x"ff"),
   949 => (x"87",x"ea",x"c0",x"49"),
   950 => (x"02",x"9b",x"4b",x"70"),
   951 => (x"8b",x"c1",x"87",x"c2"),
   952 => (x"c8",x"48",x"d0",x"ff"),
   953 => (x"d5",x"c1",x"78",x"c5"),
   954 => (x"c6",x"49",x"73",x"7c"),
   955 => (x"e7",x"e5",x"c2",x"31"),
   956 => (x"48",x"4a",x"bf",x"97"),
   957 => (x"7c",x"70",x"b0",x"71"),
   958 => (x"c4",x"48",x"d0",x"ff"),
   959 => (x"fe",x"48",x"73",x"78"),
   960 => (x"5e",x"0e",x"87",x"d5"),
   961 => (x"0e",x"5d",x"5c",x"5b"),
   962 => (x"4c",x"71",x"86",x"f4"),
   963 => (x"c0",x"48",x"a6",x"c4"),
   964 => (x"7e",x"a4",x"c8",x"78"),
   965 => (x"49",x"bf",x"97",x"6e"),
   966 => (x"05",x"a9",x"c1",x"c1"),
   967 => (x"a4",x"c9",x"87",x"dd"),
   968 => (x"49",x"69",x"97",x"49"),
   969 => (x"05",x"a9",x"d2",x"c1"),
   970 => (x"a4",x"ca",x"87",x"d1"),
   971 => (x"49",x"69",x"97",x"49"),
   972 => (x"05",x"a9",x"c3",x"c1"),
   973 => (x"48",x"df",x"87",x"c5"),
   974 => (x"fa",x"87",x"e1",x"c2"),
   975 => (x"4b",x"c0",x"87",x"e7"),
   976 => (x"97",x"e1",x"ff",x"c0"),
   977 => (x"a9",x"c0",x"49",x"bf"),
   978 => (x"fb",x"87",x"cf",x"04"),
   979 => (x"83",x"c1",x"87",x"cc"),
   980 => (x"97",x"e1",x"ff",x"c0"),
   981 => (x"06",x"ab",x"49",x"bf"),
   982 => (x"ff",x"c0",x"87",x"f1"),
   983 => (x"02",x"bf",x"97",x"e1"),
   984 => (x"e0",x"f9",x"87",x"cf"),
   985 => (x"99",x"49",x"70",x"87"),
   986 => (x"c0",x"87",x"c6",x"02"),
   987 => (x"f1",x"05",x"a9",x"ec"),
   988 => (x"f9",x"4b",x"c0",x"87"),
   989 => (x"4d",x"70",x"87",x"cf"),
   990 => (x"cc",x"87",x"ca",x"f9"),
   991 => (x"c4",x"f9",x"58",x"a6"),
   992 => (x"c1",x"4a",x"70",x"87"),
   993 => (x"bf",x"97",x"6e",x"83"),
   994 => (x"c7",x"02",x"ad",x"49"),
   995 => (x"ad",x"ff",x"c0",x"87"),
   996 => (x"87",x"ea",x"c0",x"05"),
   997 => (x"97",x"49",x"a4",x"c9"),
   998 => (x"66",x"c8",x"49",x"69"),
   999 => (x"87",x"c7",x"02",x"a9"),
  1000 => (x"a8",x"ff",x"c0",x"48"),
  1001 => (x"ca",x"87",x"d7",x"05"),
  1002 => (x"69",x"97",x"49",x"a4"),
  1003 => (x"c6",x"02",x"aa",x"49"),
  1004 => (x"aa",x"ff",x"c0",x"87"),
  1005 => (x"c4",x"87",x"c7",x"05"),
  1006 => (x"78",x"c1",x"48",x"a6"),
  1007 => (x"ec",x"c0",x"87",x"d3"),
  1008 => (x"87",x"c6",x"02",x"ad"),
  1009 => (x"05",x"ad",x"fb",x"c0"),
  1010 => (x"4b",x"c0",x"87",x"c7"),
  1011 => (x"c1",x"48",x"a6",x"c4"),
  1012 => (x"02",x"66",x"c4",x"78"),
  1013 => (x"f8",x"87",x"dc",x"fe"),
  1014 => (x"48",x"73",x"87",x"f7"),
  1015 => (x"f4",x"fa",x"8e",x"f4"),
  1016 => (x"5e",x"0e",x"00",x"87"),
  1017 => (x"0e",x"5d",x"5c",x"5b"),
  1018 => (x"c0",x"4b",x"71",x"1e"),
  1019 => (x"04",x"ab",x"4d",x"4c"),
  1020 => (x"c0",x"87",x"e8",x"c0"),
  1021 => (x"75",x"1e",x"c2",x"fc"),
  1022 => (x"87",x"c4",x"02",x"9d"),
  1023 => (x"87",x"c2",x"4a",x"c0"),
  1024 => (x"49",x"72",x"4a",x"c1"),
  1025 => (x"c4",x"87",x"c8",x"ef"),
  1026 => (x"c1",x"7e",x"70",x"86"),
  1027 => (x"c2",x"05",x"6e",x"84"),
  1028 => (x"c1",x"4c",x"73",x"87"),
  1029 => (x"06",x"ac",x"73",x"85"),
  1030 => (x"6e",x"87",x"d8",x"ff"),
  1031 => (x"4d",x"26",x"26",x"48"),
  1032 => (x"4b",x"26",x"4c",x"26"),
  1033 => (x"5e",x"0e",x"4f",x"26"),
  1034 => (x"0e",x"5d",x"5c",x"5b"),
  1035 => (x"49",x"4c",x"71",x"1e"),
  1036 => (x"c9",x"c3",x"91",x"de"),
  1037 => (x"85",x"71",x"4d",x"c1"),
  1038 => (x"c1",x"02",x"6d",x"97"),
  1039 => (x"c8",x"c3",x"87",x"dd"),
  1040 => (x"74",x"4a",x"bf",x"ec"),
  1041 => (x"fe",x"49",x"72",x"82"),
  1042 => (x"7e",x"70",x"87",x"d8"),
  1043 => (x"f3",x"c0",x"02",x"6e"),
  1044 => (x"f4",x"c8",x"c3",x"87"),
  1045 => (x"cb",x"4a",x"6e",x"4b"),
  1046 => (x"cb",x"c1",x"ff",x"49"),
  1047 => (x"cb",x"4b",x"74",x"87"),
  1048 => (x"ee",x"e2",x"c1",x"93"),
  1049 => (x"c1",x"83",x"c4",x"83"),
  1050 => (x"74",x"7b",x"df",x"c2"),
  1051 => (x"d6",x"cc",x"c1",x"49"),
  1052 => (x"c3",x"7b",x"75",x"87"),
  1053 => (x"bf",x"97",x"c0",x"c9"),
  1054 => (x"c8",x"c3",x"1e",x"49"),
  1055 => (x"e3",x"c1",x"49",x"f4"),
  1056 => (x"86",x"c4",x"87",x"d6"),
  1057 => (x"cb",x"c1",x"49",x"74"),
  1058 => (x"49",x"c0",x"87",x"fd"),
  1059 => (x"87",x"dc",x"cd",x"c1"),
  1060 => (x"48",x"e8",x"c8",x"c3"),
  1061 => (x"49",x"c1",x"78",x"c0"),
  1062 => (x"26",x"87",x"fe",x"dc"),
  1063 => (x"4c",x"87",x"ff",x"fd"),
  1064 => (x"69",x"64",x"61",x"6f"),
  1065 => (x"2e",x"2e",x"67",x"6e"),
  1066 => (x"5e",x"0e",x"00",x"2e"),
  1067 => (x"71",x"0e",x"5c",x"5b"),
  1068 => (x"c8",x"c3",x"4a",x"4b"),
  1069 => (x"72",x"82",x"bf",x"ec"),
  1070 => (x"87",x"e6",x"fc",x"49"),
  1071 => (x"02",x"9c",x"4c",x"70"),
  1072 => (x"eb",x"49",x"87",x"c4"),
  1073 => (x"c8",x"c3",x"87",x"d1"),
  1074 => (x"78",x"c0",x"48",x"ec"),
  1075 => (x"c8",x"dc",x"49",x"c1"),
  1076 => (x"87",x"cc",x"fd",x"87"),
  1077 => (x"5c",x"5b",x"5e",x"0e"),
  1078 => (x"86",x"f4",x"0e",x"5d"),
  1079 => (x"4d",x"f6",x"fb",x"c2"),
  1080 => (x"a6",x"c4",x"4c",x"c0"),
  1081 => (x"c3",x"78",x"c0",x"48"),
  1082 => (x"49",x"bf",x"ec",x"c8"),
  1083 => (x"c1",x"06",x"a9",x"c0"),
  1084 => (x"fb",x"c2",x"87",x"c1"),
  1085 => (x"02",x"98",x"48",x"f6"),
  1086 => (x"c0",x"87",x"f8",x"c0"),
  1087 => (x"c8",x"1e",x"c2",x"fc"),
  1088 => (x"87",x"c7",x"02",x"66"),
  1089 => (x"c0",x"48",x"a6",x"c4"),
  1090 => (x"c4",x"87",x"c5",x"78"),
  1091 => (x"78",x"c1",x"48",x"a6"),
  1092 => (x"ea",x"49",x"66",x"c4"),
  1093 => (x"86",x"c4",x"87",x"f9"),
  1094 => (x"84",x"c1",x"4d",x"70"),
  1095 => (x"c1",x"48",x"66",x"c4"),
  1096 => (x"58",x"a6",x"c8",x"80"),
  1097 => (x"bf",x"ec",x"c8",x"c3"),
  1098 => (x"c6",x"03",x"ac",x"49"),
  1099 => (x"05",x"9d",x"75",x"87"),
  1100 => (x"c0",x"87",x"c8",x"ff"),
  1101 => (x"02",x"9d",x"75",x"4c"),
  1102 => (x"c0",x"87",x"e0",x"c3"),
  1103 => (x"c8",x"1e",x"c2",x"fc"),
  1104 => (x"87",x"c7",x"02",x"66"),
  1105 => (x"c0",x"48",x"a6",x"cc"),
  1106 => (x"cc",x"87",x"c5",x"78"),
  1107 => (x"78",x"c1",x"48",x"a6"),
  1108 => (x"e9",x"49",x"66",x"cc"),
  1109 => (x"86",x"c4",x"87",x"f9"),
  1110 => (x"02",x"6e",x"7e",x"70"),
  1111 => (x"6e",x"87",x"e9",x"c2"),
  1112 => (x"97",x"81",x"cb",x"49"),
  1113 => (x"99",x"d0",x"49",x"69"),
  1114 => (x"87",x"d6",x"c1",x"02"),
  1115 => (x"4a",x"ea",x"c2",x"c1"),
  1116 => (x"91",x"cb",x"49",x"74"),
  1117 => (x"81",x"ee",x"e2",x"c1"),
  1118 => (x"81",x"c8",x"79",x"72"),
  1119 => (x"74",x"51",x"ff",x"c3"),
  1120 => (x"c3",x"91",x"de",x"49"),
  1121 => (x"71",x"4d",x"c1",x"c9"),
  1122 => (x"97",x"c1",x"c2",x"85"),
  1123 => (x"49",x"a5",x"c1",x"7d"),
  1124 => (x"c3",x"51",x"e0",x"c0"),
  1125 => (x"bf",x"97",x"c6",x"c4"),
  1126 => (x"c1",x"87",x"d2",x"02"),
  1127 => (x"4b",x"a5",x"c2",x"84"),
  1128 => (x"4a",x"c6",x"c4",x"c3"),
  1129 => (x"fb",x"fe",x"49",x"db"),
  1130 => (x"db",x"c1",x"87",x"fe"),
  1131 => (x"49",x"a5",x"cd",x"87"),
  1132 => (x"84",x"c1",x"51",x"c0"),
  1133 => (x"6e",x"4b",x"a5",x"c2"),
  1134 => (x"fe",x"49",x"cb",x"4a"),
  1135 => (x"c1",x"87",x"e9",x"fb"),
  1136 => (x"c0",x"c1",x"87",x"c6"),
  1137 => (x"49",x"74",x"4a",x"e6"),
  1138 => (x"e2",x"c1",x"91",x"cb"),
  1139 => (x"79",x"72",x"81",x"ee"),
  1140 => (x"97",x"c6",x"c4",x"c3"),
  1141 => (x"87",x"d8",x"02",x"bf"),
  1142 => (x"91",x"de",x"49",x"74"),
  1143 => (x"c9",x"c3",x"84",x"c1"),
  1144 => (x"83",x"71",x"4b",x"c1"),
  1145 => (x"4a",x"c6",x"c4",x"c3"),
  1146 => (x"fa",x"fe",x"49",x"dd"),
  1147 => (x"87",x"d8",x"87",x"fa"),
  1148 => (x"93",x"de",x"4b",x"74"),
  1149 => (x"83",x"c1",x"c9",x"c3"),
  1150 => (x"c0",x"49",x"a3",x"cb"),
  1151 => (x"73",x"84",x"c1",x"51"),
  1152 => (x"49",x"cb",x"4a",x"6e"),
  1153 => (x"87",x"e0",x"fa",x"fe"),
  1154 => (x"c1",x"48",x"66",x"c4"),
  1155 => (x"58",x"a6",x"c8",x"80"),
  1156 => (x"c0",x"03",x"ac",x"c7"),
  1157 => (x"05",x"6e",x"87",x"c5"),
  1158 => (x"74",x"87",x"e0",x"fc"),
  1159 => (x"f7",x"8e",x"f4",x"48"),
  1160 => (x"73",x"1e",x"87",x"fc"),
  1161 => (x"49",x"4b",x"71",x"1e"),
  1162 => (x"e2",x"c1",x"91",x"cb"),
  1163 => (x"a1",x"c8",x"81",x"ee"),
  1164 => (x"e7",x"e5",x"c2",x"4a"),
  1165 => (x"c9",x"50",x"12",x"48"),
  1166 => (x"ff",x"c0",x"4a",x"a1"),
  1167 => (x"50",x"12",x"48",x"e1"),
  1168 => (x"c9",x"c3",x"81",x"ca"),
  1169 => (x"50",x"11",x"48",x"c0"),
  1170 => (x"97",x"c0",x"c9",x"c3"),
  1171 => (x"c0",x"1e",x"49",x"bf"),
  1172 => (x"c3",x"dc",x"c1",x"49"),
  1173 => (x"e8",x"c8",x"c3",x"87"),
  1174 => (x"c1",x"78",x"de",x"48"),
  1175 => (x"87",x"f9",x"d5",x"49"),
  1176 => (x"87",x"fe",x"f6",x"26"),
  1177 => (x"49",x"4a",x"71",x"1e"),
  1178 => (x"e2",x"c1",x"91",x"cb"),
  1179 => (x"81",x"c8",x"81",x"ee"),
  1180 => (x"c8",x"c3",x"48",x"11"),
  1181 => (x"c8",x"c3",x"58",x"ec"),
  1182 => (x"78",x"c0",x"48",x"ec"),
  1183 => (x"d8",x"d5",x"49",x"c1"),
  1184 => (x"1e",x"4f",x"26",x"87"),
  1185 => (x"c5",x"c1",x"49",x"c0"),
  1186 => (x"4f",x"26",x"87",x"e2"),
  1187 => (x"02",x"99",x"71",x"1e"),
  1188 => (x"e4",x"c1",x"87",x"d2"),
  1189 => (x"50",x"c0",x"48",x"c3"),
  1190 => (x"c9",x"c1",x"80",x"f7"),
  1191 => (x"e2",x"c1",x"40",x"e4"),
  1192 => (x"87",x"ce",x"78",x"e7"),
  1193 => (x"48",x"ff",x"e3",x"c1"),
  1194 => (x"78",x"e0",x"e2",x"c1"),
  1195 => (x"ca",x"c1",x"80",x"fc"),
  1196 => (x"4f",x"26",x"78",x"c3"),
  1197 => (x"5c",x"5b",x"5e",x"0e"),
  1198 => (x"4a",x"4c",x"71",x"0e"),
  1199 => (x"e2",x"c1",x"92",x"cb"),
  1200 => (x"a2",x"c8",x"82",x"ee"),
  1201 => (x"4b",x"a2",x"c9",x"49"),
  1202 => (x"1e",x"4b",x"6b",x"97"),
  1203 => (x"1e",x"49",x"69",x"97"),
  1204 => (x"49",x"12",x"82",x"ca"),
  1205 => (x"87",x"c3",x"e6",x"c0"),
  1206 => (x"fc",x"d3",x"49",x"c0"),
  1207 => (x"c1",x"49",x"74",x"87"),
  1208 => (x"f8",x"87",x"e4",x"c2"),
  1209 => (x"87",x"f8",x"f4",x"8e"),
  1210 => (x"71",x"1e",x"73",x"1e"),
  1211 => (x"4a",x"a3",x"c6",x"4b"),
  1212 => (x"c1",x"87",x"db",x"02"),
  1213 => (x"87",x"d6",x"02",x"8a"),
  1214 => (x"da",x"c1",x"02",x"8a"),
  1215 => (x"c0",x"02",x"8a",x"87"),
  1216 => (x"02",x"8a",x"87",x"fc"),
  1217 => (x"8a",x"87",x"e1",x"c0"),
  1218 => (x"c1",x"87",x"cb",x"02"),
  1219 => (x"49",x"c7",x"87",x"db"),
  1220 => (x"c1",x"87",x"d1",x"fd"),
  1221 => (x"c8",x"c3",x"87",x"de"),
  1222 => (x"c1",x"02",x"bf",x"ec"),
  1223 => (x"c1",x"48",x"87",x"cb"),
  1224 => (x"f0",x"c8",x"c3",x"88"),
  1225 => (x"87",x"c1",x"c1",x"58"),
  1226 => (x"bf",x"f0",x"c8",x"c3"),
  1227 => (x"87",x"f9",x"c0",x"02"),
  1228 => (x"bf",x"ec",x"c8",x"c3"),
  1229 => (x"c3",x"80",x"c1",x"48"),
  1230 => (x"c0",x"58",x"f0",x"c8"),
  1231 => (x"c8",x"c3",x"87",x"eb"),
  1232 => (x"c6",x"49",x"bf",x"ec"),
  1233 => (x"f0",x"c8",x"c3",x"89"),
  1234 => (x"a9",x"b7",x"c0",x"59"),
  1235 => (x"c3",x"87",x"da",x"03"),
  1236 => (x"c0",x"48",x"ec",x"c8"),
  1237 => (x"c3",x"87",x"d2",x"78"),
  1238 => (x"02",x"bf",x"f0",x"c8"),
  1239 => (x"c8",x"c3",x"87",x"cb"),
  1240 => (x"c6",x"48",x"bf",x"ec"),
  1241 => (x"f0",x"c8",x"c3",x"80"),
  1242 => (x"d1",x"49",x"c0",x"58"),
  1243 => (x"49",x"73",x"87",x"eb"),
  1244 => (x"87",x"d3",x"c0",x"c1"),
  1245 => (x"1e",x"87",x"eb",x"f2"),
  1246 => (x"4b",x"71",x"1e",x"73"),
  1247 => (x"48",x"e8",x"c8",x"c3"),
  1248 => (x"49",x"c0",x"78",x"dd"),
  1249 => (x"73",x"87",x"d2",x"d1"),
  1250 => (x"fa",x"ff",x"c0",x"49"),
  1251 => (x"87",x"d2",x"f2",x"87"),
  1252 => (x"5c",x"5b",x"5e",x"0e"),
  1253 => (x"cc",x"4c",x"71",x"0e"),
  1254 => (x"4b",x"74",x"1e",x"66"),
  1255 => (x"e2",x"c1",x"93",x"cb"),
  1256 => (x"a3",x"c4",x"83",x"ee"),
  1257 => (x"fe",x"49",x"6a",x"4a"),
  1258 => (x"c1",x"87",x"cd",x"f4"),
  1259 => (x"c8",x"7b",x"e2",x"c8"),
  1260 => (x"66",x"d4",x"49",x"a3"),
  1261 => (x"49",x"a3",x"c9",x"51"),
  1262 => (x"ca",x"51",x"66",x"d8"),
  1263 => (x"66",x"dc",x"49",x"a3"),
  1264 => (x"db",x"f1",x"26",x"51"),
  1265 => (x"5b",x"5e",x"0e",x"87"),
  1266 => (x"ff",x"0e",x"5d",x"5c"),
  1267 => (x"a6",x"dc",x"86",x"cc"),
  1268 => (x"48",x"a6",x"c8",x"59"),
  1269 => (x"80",x"c4",x"78",x"c0"),
  1270 => (x"78",x"66",x"c8",x"c1"),
  1271 => (x"78",x"c1",x"80",x"c4"),
  1272 => (x"78",x"c1",x"80",x"c4"),
  1273 => (x"48",x"f0",x"c8",x"c3"),
  1274 => (x"c8",x"c3",x"78",x"c1"),
  1275 => (x"de",x"48",x"bf",x"e8"),
  1276 => (x"87",x"cb",x"05",x"a8"),
  1277 => (x"70",x"87",x"dd",x"f3"),
  1278 => (x"59",x"a6",x"cc",x"49"),
  1279 => (x"e7",x"87",x"d6",x"ce"),
  1280 => (x"d5",x"e8",x"87",x"e3"),
  1281 => (x"87",x"fd",x"e6",x"87"),
  1282 => (x"fb",x"c0",x"4c",x"70"),
  1283 => (x"d8",x"c1",x"02",x"ac"),
  1284 => (x"05",x"66",x"d8",x"87"),
  1285 => (x"c0",x"87",x"ca",x"c1"),
  1286 => (x"1e",x"c1",x"1e",x"1e"),
  1287 => (x"1e",x"d1",x"e4",x"c1"),
  1288 => (x"eb",x"fd",x"49",x"c0"),
  1289 => (x"c0",x"86",x"d0",x"87"),
  1290 => (x"d9",x"02",x"ac",x"fb"),
  1291 => (x"66",x"c4",x"c1",x"87"),
  1292 => (x"6a",x"82",x"c4",x"4a"),
  1293 => (x"74",x"81",x"c7",x"49"),
  1294 => (x"d8",x"1e",x"c1",x"51"),
  1295 => (x"c8",x"49",x"6a",x"1e"),
  1296 => (x"87",x"ea",x"e7",x"81"),
  1297 => (x"c8",x"c1",x"86",x"c8"),
  1298 => (x"a8",x"c0",x"48",x"66"),
  1299 => (x"c8",x"87",x"c7",x"01"),
  1300 => (x"78",x"c1",x"48",x"a6"),
  1301 => (x"c8",x"c1",x"87",x"ce"),
  1302 => (x"88",x"c1",x"48",x"66"),
  1303 => (x"c3",x"58",x"a6",x"d0"),
  1304 => (x"87",x"f6",x"e6",x"87"),
  1305 => (x"c2",x"48",x"a6",x"d0"),
  1306 => (x"02",x"9c",x"74",x"78"),
  1307 => (x"c8",x"87",x"e2",x"cc"),
  1308 => (x"cc",x"c1",x"48",x"66"),
  1309 => (x"cc",x"03",x"a8",x"66"),
  1310 => (x"a6",x"dc",x"87",x"d7"),
  1311 => (x"e5",x"78",x"c0",x"48"),
  1312 => (x"4c",x"70",x"87",x"c3"),
  1313 => (x"dd",x"48",x"66",x"d8"),
  1314 => (x"87",x"c6",x"05",x"a8"),
  1315 => (x"d8",x"48",x"a6",x"dc"),
  1316 => (x"d0",x"c1",x"78",x"66"),
  1317 => (x"e8",x"c0",x"05",x"ac"),
  1318 => (x"87",x"e9",x"e4",x"87"),
  1319 => (x"70",x"87",x"e6",x"e4"),
  1320 => (x"ac",x"ec",x"c0",x"4c"),
  1321 => (x"e5",x"87",x"c5",x"05"),
  1322 => (x"4c",x"70",x"87",x"f0"),
  1323 => (x"05",x"ac",x"d0",x"c1"),
  1324 => (x"66",x"d4",x"87",x"c8"),
  1325 => (x"d8",x"80",x"c1",x"48"),
  1326 => (x"d0",x"c1",x"58",x"a6"),
  1327 => (x"d8",x"ff",x"02",x"ac"),
  1328 => (x"a6",x"e0",x"c0",x"87"),
  1329 => (x"78",x"66",x"d8",x"48"),
  1330 => (x"c0",x"48",x"66",x"dc"),
  1331 => (x"05",x"a8",x"66",x"e0"),
  1332 => (x"c4",x"87",x"d0",x"ca"),
  1333 => (x"f0",x"c0",x"48",x"a6"),
  1334 => (x"80",x"e0",x"c0",x"78"),
  1335 => (x"c4",x"78",x"66",x"d0"),
  1336 => (x"c4",x"78",x"c0",x"80"),
  1337 => (x"74",x"78",x"c0",x"80"),
  1338 => (x"8d",x"fb",x"c0",x"4d"),
  1339 => (x"87",x"cc",x"c9",x"02"),
  1340 => (x"db",x"02",x"8d",x"c9"),
  1341 => (x"02",x"8d",x"c2",x"87"),
  1342 => (x"c9",x"87",x"cd",x"c1"),
  1343 => (x"d1",x"c4",x"02",x"8d"),
  1344 => (x"02",x"8d",x"c4",x"87"),
  1345 => (x"c1",x"87",x"c6",x"c1"),
  1346 => (x"c5",x"c4",x"02",x"8d"),
  1347 => (x"87",x"e6",x"c8",x"87"),
  1348 => (x"cb",x"49",x"66",x"c8"),
  1349 => (x"66",x"c4",x"c1",x"91"),
  1350 => (x"4a",x"a1",x"c4",x"81"),
  1351 => (x"1e",x"71",x"7e",x"6a"),
  1352 => (x"48",x"cc",x"df",x"c1"),
  1353 => (x"cc",x"49",x"66",x"c4"),
  1354 => (x"41",x"20",x"4a",x"a1"),
  1355 => (x"ff",x"05",x"aa",x"71"),
  1356 => (x"51",x"10",x"87",x"f8"),
  1357 => (x"cd",x"c1",x"49",x"26"),
  1358 => (x"dd",x"e3",x"79",x"f7"),
  1359 => (x"c0",x"4c",x"70",x"87"),
  1360 => (x"c1",x"48",x"a6",x"ec"),
  1361 => (x"87",x"f4",x"c7",x"78"),
  1362 => (x"c0",x"48",x"a6",x"c4"),
  1363 => (x"48",x"66",x"d0",x"78"),
  1364 => (x"a6",x"d4",x"80",x"c1"),
  1365 => (x"87",x"ed",x"e1",x"58"),
  1366 => (x"ec",x"c0",x"4c",x"70"),
  1367 => (x"87",x"d4",x"02",x"ac"),
  1368 => (x"c0",x"02",x"66",x"c4"),
  1369 => (x"a6",x"c8",x"87",x"c5"),
  1370 => (x"74",x"87",x"c9",x"5c"),
  1371 => (x"88",x"f0",x"c0",x"48"),
  1372 => (x"58",x"a6",x"e8",x"c0"),
  1373 => (x"02",x"ac",x"ec",x"c0"),
  1374 => (x"c8",x"e1",x"87",x"cc"),
  1375 => (x"c0",x"4c",x"70",x"87"),
  1376 => (x"ff",x"05",x"ac",x"ec"),
  1377 => (x"66",x"c4",x"87",x"f4"),
  1378 => (x"49",x"66",x"d8",x"1e"),
  1379 => (x"66",x"ec",x"c0",x"1e"),
  1380 => (x"d1",x"e4",x"c1",x"1e"),
  1381 => (x"49",x"66",x"d8",x"1e"),
  1382 => (x"c0",x"87",x"f5",x"f7"),
  1383 => (x"c0",x"1e",x"ca",x"1e"),
  1384 => (x"cb",x"49",x"66",x"e0"),
  1385 => (x"66",x"dc",x"c1",x"91"),
  1386 => (x"48",x"a6",x"d8",x"81"),
  1387 => (x"d8",x"78",x"a1",x"c4"),
  1388 => (x"e1",x"49",x"bf",x"66"),
  1389 => (x"86",x"d8",x"87",x"f8"),
  1390 => (x"06",x"a8",x"b7",x"c0"),
  1391 => (x"c1",x"87",x"ca",x"c1"),
  1392 => (x"c8",x"1e",x"de",x"1e"),
  1393 => (x"e1",x"49",x"bf",x"66"),
  1394 => (x"86",x"c8",x"87",x"e4"),
  1395 => (x"c0",x"48",x"49",x"70"),
  1396 => (x"e8",x"c0",x"88",x"08"),
  1397 => (x"b7",x"c0",x"58",x"a6"),
  1398 => (x"ec",x"c0",x"06",x"a8"),
  1399 => (x"66",x"e4",x"c0",x"87"),
  1400 => (x"a8",x"b7",x"dd",x"48"),
  1401 => (x"87",x"e1",x"c0",x"03"),
  1402 => (x"c0",x"49",x"bf",x"6e"),
  1403 => (x"c0",x"81",x"66",x"e4"),
  1404 => (x"e4",x"c0",x"51",x"e0"),
  1405 => (x"81",x"c1",x"49",x"66"),
  1406 => (x"c2",x"81",x"bf",x"6e"),
  1407 => (x"e4",x"c0",x"51",x"c1"),
  1408 => (x"81",x"c2",x"49",x"66"),
  1409 => (x"c0",x"81",x"bf",x"6e"),
  1410 => (x"a6",x"ec",x"c0",x"51"),
  1411 => (x"c4",x"78",x"c1",x"48"),
  1412 => (x"c8",x"e2",x"87",x"ea"),
  1413 => (x"a6",x"e8",x"c0",x"87"),
  1414 => (x"87",x"c1",x"e2",x"58"),
  1415 => (x"58",x"a6",x"f0",x"c0"),
  1416 => (x"05",x"a8",x"ec",x"c0"),
  1417 => (x"a6",x"87",x"c9",x"c0"),
  1418 => (x"66",x"e4",x"c0",x"48"),
  1419 => (x"87",x"c4",x"c0",x"78"),
  1420 => (x"87",x"d1",x"de",x"ff"),
  1421 => (x"cb",x"49",x"66",x"c8"),
  1422 => (x"66",x"c4",x"c1",x"91"),
  1423 => (x"c8",x"80",x"71",x"48"),
  1424 => (x"66",x"c4",x"58",x"a6"),
  1425 => (x"c4",x"82",x"c8",x"4a"),
  1426 => (x"81",x"ca",x"49",x"66"),
  1427 => (x"51",x"66",x"e4",x"c0"),
  1428 => (x"49",x"66",x"ec",x"c0"),
  1429 => (x"e4",x"c0",x"81",x"c1"),
  1430 => (x"48",x"c1",x"89",x"66"),
  1431 => (x"49",x"70",x"30",x"71"),
  1432 => (x"97",x"71",x"89",x"c1"),
  1433 => (x"dd",x"cc",x"c3",x"7a"),
  1434 => (x"e4",x"c0",x"49",x"bf"),
  1435 => (x"6a",x"97",x"29",x"66"),
  1436 => (x"98",x"71",x"48",x"4a"),
  1437 => (x"58",x"a6",x"f4",x"c0"),
  1438 => (x"c4",x"49",x"66",x"c4"),
  1439 => (x"c0",x"7e",x"69",x"81"),
  1440 => (x"dc",x"48",x"66",x"e0"),
  1441 => (x"c0",x"02",x"a8",x"66"),
  1442 => (x"a6",x"dc",x"87",x"c8"),
  1443 => (x"c0",x"78",x"c0",x"48"),
  1444 => (x"a6",x"dc",x"87",x"c5"),
  1445 => (x"dc",x"78",x"c1",x"48"),
  1446 => (x"e0",x"c0",x"1e",x"66"),
  1447 => (x"49",x"66",x"c8",x"1e"),
  1448 => (x"87",x"ca",x"de",x"ff"),
  1449 => (x"4c",x"70",x"86",x"c8"),
  1450 => (x"06",x"ac",x"b7",x"c0"),
  1451 => (x"6e",x"87",x"d6",x"c1"),
  1452 => (x"70",x"80",x"74",x"48"),
  1453 => (x"49",x"e0",x"c0",x"7e"),
  1454 => (x"4b",x"6e",x"89",x"74"),
  1455 => (x"4a",x"c9",x"df",x"c1"),
  1456 => (x"e3",x"e7",x"fe",x"71"),
  1457 => (x"c2",x"48",x"6e",x"87"),
  1458 => (x"c0",x"7e",x"70",x"80"),
  1459 => (x"c1",x"48",x"66",x"e8"),
  1460 => (x"a6",x"ec",x"c0",x"80"),
  1461 => (x"66",x"f0",x"c0",x"58"),
  1462 => (x"70",x"81",x"c1",x"49"),
  1463 => (x"c5",x"c0",x"02",x"a9"),
  1464 => (x"c0",x"4d",x"c0",x"87"),
  1465 => (x"4d",x"c1",x"87",x"c2"),
  1466 => (x"a4",x"c2",x"1e",x"75"),
  1467 => (x"48",x"e0",x"c0",x"49"),
  1468 => (x"49",x"70",x"88",x"71"),
  1469 => (x"49",x"66",x"c8",x"1e"),
  1470 => (x"87",x"f2",x"dc",x"ff"),
  1471 => (x"b7",x"c0",x"86",x"c8"),
  1472 => (x"c6",x"ff",x"01",x"a8"),
  1473 => (x"66",x"e8",x"c0",x"87"),
  1474 => (x"87",x"d3",x"c0",x"02"),
  1475 => (x"c9",x"49",x"66",x"c4"),
  1476 => (x"66",x"e8",x"c0",x"81"),
  1477 => (x"48",x"66",x"c4",x"51"),
  1478 => (x"78",x"f4",x"ca",x"c1"),
  1479 => (x"c4",x"87",x"ce",x"c0"),
  1480 => (x"81",x"c9",x"49",x"66"),
  1481 => (x"66",x"c4",x"51",x"c2"),
  1482 => (x"ce",x"f5",x"c2",x"48"),
  1483 => (x"a6",x"ec",x"c0",x"78"),
  1484 => (x"c0",x"78",x"c1",x"48"),
  1485 => (x"db",x"ff",x"87",x"c6"),
  1486 => (x"4c",x"70",x"87",x"e0"),
  1487 => (x"02",x"66",x"ec",x"c0"),
  1488 => (x"c8",x"87",x"f5",x"c0"),
  1489 => (x"66",x"cc",x"48",x"66"),
  1490 => (x"cb",x"c0",x"04",x"a8"),
  1491 => (x"48",x"66",x"c8",x"87"),
  1492 => (x"a6",x"cc",x"80",x"c1"),
  1493 => (x"87",x"e0",x"c0",x"58"),
  1494 => (x"c1",x"48",x"66",x"cc"),
  1495 => (x"58",x"a6",x"d0",x"88"),
  1496 => (x"c1",x"87",x"d5",x"c0"),
  1497 => (x"c0",x"05",x"ac",x"c6"),
  1498 => (x"66",x"d0",x"87",x"c8"),
  1499 => (x"d4",x"80",x"c1",x"48"),
  1500 => (x"da",x"ff",x"58",x"a6"),
  1501 => (x"4c",x"70",x"87",x"e4"),
  1502 => (x"c1",x"48",x"66",x"d4"),
  1503 => (x"58",x"a6",x"d8",x"80"),
  1504 => (x"c0",x"02",x"9c",x"74"),
  1505 => (x"66",x"c8",x"87",x"cb"),
  1506 => (x"66",x"cc",x"c1",x"48"),
  1507 => (x"e9",x"f3",x"04",x"a8"),
  1508 => (x"fc",x"d9",x"ff",x"87"),
  1509 => (x"48",x"66",x"c8",x"87"),
  1510 => (x"c0",x"03",x"a8",x"c7"),
  1511 => (x"c8",x"c3",x"87",x"e5"),
  1512 => (x"78",x"c0",x"48",x"f0"),
  1513 => (x"cb",x"49",x"66",x"c8"),
  1514 => (x"66",x"c4",x"c1",x"91"),
  1515 => (x"4a",x"a1",x"c4",x"81"),
  1516 => (x"52",x"c0",x"4a",x"6a"),
  1517 => (x"48",x"66",x"c8",x"79"),
  1518 => (x"a6",x"cc",x"80",x"c1"),
  1519 => (x"04",x"a8",x"c7",x"58"),
  1520 => (x"ff",x"87",x"db",x"ff"),
  1521 => (x"d5",x"e1",x"8e",x"cc"),
  1522 => (x"00",x"20",x"3a",x"87"),
  1523 => (x"20",x"50",x"49",x"44"),
  1524 => (x"74",x"69",x"77",x"53"),
  1525 => (x"73",x"65",x"68",x"63"),
  1526 => (x"1e",x"73",x"1e",x"00"),
  1527 => (x"02",x"9b",x"4b",x"71"),
  1528 => (x"c8",x"c3",x"87",x"c6"),
  1529 => (x"78",x"c0",x"48",x"ec"),
  1530 => (x"c8",x"c3",x"1e",x"c7"),
  1531 => (x"1e",x"49",x"bf",x"ec"),
  1532 => (x"1e",x"ee",x"e2",x"c1"),
  1533 => (x"bf",x"e8",x"c8",x"c3"),
  1534 => (x"87",x"c9",x"ef",x"49"),
  1535 => (x"c8",x"c3",x"86",x"cc"),
  1536 => (x"ea",x"49",x"bf",x"e8"),
  1537 => (x"9b",x"73",x"87",x"c6"),
  1538 => (x"c1",x"87",x"c8",x"02"),
  1539 => (x"c0",x"49",x"ee",x"e2"),
  1540 => (x"e0",x"87",x"c6",x"ef"),
  1541 => (x"c7",x"1e",x"87",x"cc"),
  1542 => (x"49",x"c1",x"87",x"d6"),
  1543 => (x"fe",x"87",x"fa",x"fe"),
  1544 => (x"70",x"87",x"f4",x"eb"),
  1545 => (x"87",x"cd",x"02",x"98"),
  1546 => (x"87",x"cf",x"f3",x"fe"),
  1547 => (x"c4",x"02",x"98",x"70"),
  1548 => (x"c2",x"4a",x"c1",x"87"),
  1549 => (x"72",x"4a",x"c0",x"87"),
  1550 => (x"87",x"ce",x"05",x"9a"),
  1551 => (x"e1",x"c1",x"1e",x"c0"),
  1552 => (x"fd",x"c0",x"49",x"eb"),
  1553 => (x"86",x"c4",x"87",x"d2"),
  1554 => (x"c5",x"c1",x"87",x"fe"),
  1555 => (x"1e",x"c0",x"87",x"c3"),
  1556 => (x"49",x"f6",x"e1",x"c1"),
  1557 => (x"87",x"c0",x"fd",x"c0"),
  1558 => (x"d4",x"c1",x"1e",x"c0"),
  1559 => (x"49",x"70",x"87",x"e8"),
  1560 => (x"87",x"f4",x"fc",x"c0"),
  1561 => (x"f8",x"87",x"c8",x"c3"),
  1562 => (x"53",x"4f",x"26",x"8e"),
  1563 => (x"61",x"66",x"20",x"44"),
  1564 => (x"64",x"65",x"6c",x"69"),
  1565 => (x"6f",x"42",x"00",x"2e"),
  1566 => (x"6e",x"69",x"74",x"6f"),
  1567 => (x"2e",x"2e",x"2e",x"67"),
  1568 => (x"f1",x"c0",x"1e",x"00"),
  1569 => (x"87",x"fa",x"87",x"fb"),
  1570 => (x"c3",x"1e",x"4f",x"26"),
  1571 => (x"c0",x"48",x"ec",x"c8"),
  1572 => (x"e8",x"c8",x"c3",x"78"),
  1573 => (x"fd",x"78",x"c0",x"48"),
  1574 => (x"87",x"e5",x"87",x"fc"),
  1575 => (x"4f",x"26",x"48",x"c0"),
  1576 => (x"78",x"45",x"20",x"80"),
  1577 => (x"80",x"00",x"74",x"69"),
  1578 => (x"63",x"61",x"42",x"20"),
  1579 => (x"12",x"64",x"00",x"6b"),
  1580 => (x"32",x"41",x"00",x"00"),
  1581 => (x"00",x"00",x"00",x"00"),
  1582 => (x"00",x"12",x"64",x"00"),
  1583 => (x"00",x"32",x"5f",x"00"),
  1584 => (x"00",x"00",x"00",x"00"),
  1585 => (x"00",x"00",x"12",x"64"),
  1586 => (x"00",x"00",x"32",x"7d"),
  1587 => (x"64",x"00",x"00",x"00"),
  1588 => (x"9b",x"00",x"00",x"12"),
  1589 => (x"00",x"00",x"00",x"32"),
  1590 => (x"12",x"64",x"00",x"00"),
  1591 => (x"32",x"b9",x"00",x"00"),
  1592 => (x"00",x"00",x"00",x"00"),
  1593 => (x"00",x"12",x"64",x"00"),
  1594 => (x"00",x"32",x"d7",x"00"),
  1595 => (x"00",x"00",x"00",x"00"),
  1596 => (x"00",x"00",x"12",x"64"),
  1597 => (x"00",x"00",x"32",x"f5"),
  1598 => (x"64",x"00",x"00",x"00"),
  1599 => (x"00",x"00",x"00",x"12"),
  1600 => (x"00",x"00",x"00",x"00"),
  1601 => (x"12",x"e8",x"00",x"00"),
  1602 => (x"00",x"00",x"00",x"00"),
  1603 => (x"00",x"00",x"00",x"00"),
  1604 => (x"61",x"6f",x"4c",x"00"),
  1605 => (x"2e",x"2a",x"20",x"64"),
  1606 => (x"f0",x"fe",x"1e",x"00"),
  1607 => (x"cd",x"78",x"c0",x"48"),
  1608 => (x"26",x"09",x"79",x"09"),
  1609 => (x"fe",x"1e",x"1e",x"4f"),
  1610 => (x"48",x"7e",x"bf",x"f0"),
  1611 => (x"1e",x"4f",x"26",x"26"),
  1612 => (x"c1",x"48",x"f0",x"fe"),
  1613 => (x"1e",x"4f",x"26",x"78"),
  1614 => (x"c0",x"48",x"f0",x"fe"),
  1615 => (x"1e",x"4f",x"26",x"78"),
  1616 => (x"52",x"c0",x"4a",x"71"),
  1617 => (x"0e",x"4f",x"26",x"52"),
  1618 => (x"5d",x"5c",x"5b",x"5e"),
  1619 => (x"71",x"86",x"f4",x"0e"),
  1620 => (x"7e",x"6d",x"97",x"4d"),
  1621 => (x"97",x"4c",x"a5",x"c1"),
  1622 => (x"a6",x"c8",x"48",x"6c"),
  1623 => (x"c4",x"48",x"6e",x"58"),
  1624 => (x"c5",x"05",x"a8",x"66"),
  1625 => (x"c0",x"48",x"ff",x"87"),
  1626 => (x"ca",x"ff",x"87",x"e6"),
  1627 => (x"49",x"a5",x"c2",x"87"),
  1628 => (x"71",x"4b",x"6c",x"97"),
  1629 => (x"6b",x"97",x"4b",x"a3"),
  1630 => (x"7e",x"6c",x"97",x"4b"),
  1631 => (x"80",x"c1",x"48",x"6e"),
  1632 => (x"c7",x"58",x"a6",x"c8"),
  1633 => (x"58",x"a6",x"cc",x"98"),
  1634 => (x"fe",x"7c",x"97",x"70"),
  1635 => (x"48",x"73",x"87",x"e1"),
  1636 => (x"4d",x"26",x"8e",x"f4"),
  1637 => (x"4b",x"26",x"4c",x"26"),
  1638 => (x"5e",x"0e",x"4f",x"26"),
  1639 => (x"f4",x"0e",x"5c",x"5b"),
  1640 => (x"d8",x"4c",x"71",x"86"),
  1641 => (x"ff",x"c3",x"4a",x"66"),
  1642 => (x"4b",x"a4",x"c2",x"9a"),
  1643 => (x"73",x"49",x"6c",x"97"),
  1644 => (x"51",x"72",x"49",x"a1"),
  1645 => (x"6e",x"7e",x"6c",x"97"),
  1646 => (x"c8",x"80",x"c1",x"48"),
  1647 => (x"98",x"c7",x"58",x"a6"),
  1648 => (x"70",x"58",x"a6",x"cc"),
  1649 => (x"ff",x"8e",x"f4",x"54"),
  1650 => (x"1e",x"1e",x"87",x"ca"),
  1651 => (x"e0",x"87",x"e8",x"fd"),
  1652 => (x"c0",x"49",x"4a",x"bf"),
  1653 => (x"02",x"99",x"c0",x"e0"),
  1654 => (x"1e",x"72",x"87",x"cb"),
  1655 => (x"49",x"d3",x"cc",x"c3"),
  1656 => (x"c4",x"87",x"f7",x"fe"),
  1657 => (x"87",x"fd",x"fc",x"86"),
  1658 => (x"c2",x"fd",x"7e",x"70"),
  1659 => (x"4f",x"26",x"26",x"87"),
  1660 => (x"d3",x"cc",x"c3",x"1e"),
  1661 => (x"87",x"c7",x"fd",x"49"),
  1662 => (x"49",x"ca",x"e7",x"c1"),
  1663 => (x"c5",x"87",x"da",x"fc"),
  1664 => (x"4f",x"26",x"87",x"d0"),
  1665 => (x"5c",x"5b",x"5e",x"0e"),
  1666 => (x"cd",x"c3",x"0e",x"5d"),
  1667 => (x"c1",x"4a",x"bf",x"e6"),
  1668 => (x"49",x"bf",x"d8",x"e9"),
  1669 => (x"71",x"bc",x"72",x"4c"),
  1670 => (x"87",x"db",x"fc",x"4d"),
  1671 => (x"49",x"74",x"4b",x"c0"),
  1672 => (x"d5",x"02",x"99",x"d0"),
  1673 => (x"d0",x"49",x"75",x"87"),
  1674 => (x"c0",x"1e",x"71",x"99"),
  1675 => (x"e1",x"ef",x"c1",x"1e"),
  1676 => (x"12",x"82",x"73",x"4a"),
  1677 => (x"87",x"e4",x"c0",x"49"),
  1678 => (x"2c",x"c1",x"86",x"c8"),
  1679 => (x"ab",x"c8",x"83",x"2d"),
  1680 => (x"87",x"da",x"ff",x"04"),
  1681 => (x"c1",x"87",x"e8",x"fb"),
  1682 => (x"c3",x"48",x"d8",x"e9"),
  1683 => (x"78",x"bf",x"e6",x"cd"),
  1684 => (x"4c",x"26",x"4d",x"26"),
  1685 => (x"4f",x"26",x"4b",x"26"),
  1686 => (x"00",x"00",x"00",x"00"),
  1687 => (x"48",x"d0",x"ff",x"1e"),
  1688 => (x"ff",x"78",x"e1",x"c8"),
  1689 => (x"78",x"c5",x"48",x"d4"),
  1690 => (x"c3",x"02",x"66",x"c4"),
  1691 => (x"78",x"e0",x"c3",x"87"),
  1692 => (x"c6",x"02",x"66",x"c8"),
  1693 => (x"48",x"d4",x"ff",x"87"),
  1694 => (x"ff",x"78",x"f0",x"c3"),
  1695 => (x"78",x"71",x"48",x"d4"),
  1696 => (x"c8",x"48",x"d0",x"ff"),
  1697 => (x"e0",x"c0",x"78",x"e1"),
  1698 => (x"0e",x"4f",x"26",x"78"),
  1699 => (x"0e",x"5c",x"5b",x"5e"),
  1700 => (x"cc",x"c3",x"4c",x"71"),
  1701 => (x"ee",x"fa",x"49",x"d3"),
  1702 => (x"c0",x"4a",x"70",x"87"),
  1703 => (x"c2",x"04",x"aa",x"b7"),
  1704 => (x"e0",x"c3",x"87",x"e3"),
  1705 => (x"87",x"c9",x"05",x"aa"),
  1706 => (x"48",x"ce",x"ed",x"c1"),
  1707 => (x"d4",x"c2",x"78",x"c1"),
  1708 => (x"aa",x"f0",x"c3",x"87"),
  1709 => (x"c1",x"87",x"c9",x"05"),
  1710 => (x"c1",x"48",x"ca",x"ed"),
  1711 => (x"87",x"f5",x"c1",x"78"),
  1712 => (x"bf",x"ce",x"ed",x"c1"),
  1713 => (x"72",x"87",x"c7",x"02"),
  1714 => (x"b3",x"c0",x"c2",x"4b"),
  1715 => (x"4b",x"72",x"87",x"c2"),
  1716 => (x"d1",x"05",x"9c",x"74"),
  1717 => (x"ca",x"ed",x"c1",x"87"),
  1718 => (x"ed",x"c1",x"1e",x"bf"),
  1719 => (x"72",x"1e",x"bf",x"ce"),
  1720 => (x"87",x"f8",x"fd",x"49"),
  1721 => (x"ed",x"c1",x"86",x"c8"),
  1722 => (x"c0",x"02",x"bf",x"ca"),
  1723 => (x"49",x"73",x"87",x"e0"),
  1724 => (x"91",x"29",x"b7",x"c4"),
  1725 => (x"81",x"e1",x"ee",x"c1"),
  1726 => (x"9a",x"cf",x"4a",x"73"),
  1727 => (x"48",x"c1",x"92",x"c2"),
  1728 => (x"4a",x"70",x"30",x"72"),
  1729 => (x"48",x"72",x"ba",x"ff"),
  1730 => (x"79",x"70",x"98",x"69"),
  1731 => (x"49",x"73",x"87",x"db"),
  1732 => (x"91",x"29",x"b7",x"c4"),
  1733 => (x"81",x"e1",x"ee",x"c1"),
  1734 => (x"9a",x"cf",x"4a",x"73"),
  1735 => (x"48",x"c3",x"92",x"c2"),
  1736 => (x"4a",x"70",x"30",x"72"),
  1737 => (x"70",x"b0",x"69",x"48"),
  1738 => (x"ce",x"ed",x"c1",x"79"),
  1739 => (x"c1",x"78",x"c0",x"48"),
  1740 => (x"c0",x"48",x"ca",x"ed"),
  1741 => (x"d3",x"cc",x"c3",x"78"),
  1742 => (x"87",x"cb",x"f8",x"49"),
  1743 => (x"b7",x"c0",x"4a",x"70"),
  1744 => (x"dd",x"fd",x"03",x"aa"),
  1745 => (x"fc",x"48",x"c0",x"87"),
  1746 => (x"00",x"00",x"87",x"c8"),
  1747 => (x"00",x"00",x"00",x"00"),
  1748 => (x"c0",x"1e",x"00",x"00"),
  1749 => (x"c4",x"49",x"72",x"4a"),
  1750 => (x"e1",x"ee",x"c1",x"91"),
  1751 => (x"c1",x"79",x"c0",x"81"),
  1752 => (x"aa",x"b7",x"d0",x"82"),
  1753 => (x"26",x"87",x"ee",x"04"),
  1754 => (x"5b",x"5e",x"0e",x"4f"),
  1755 => (x"71",x"0e",x"5d",x"5c"),
  1756 => (x"87",x"c3",x"f7",x"4d"),
  1757 => (x"b7",x"c4",x"4a",x"75"),
  1758 => (x"ee",x"c1",x"92",x"2a"),
  1759 => (x"4c",x"75",x"82",x"e1"),
  1760 => (x"94",x"c2",x"9c",x"cf"),
  1761 => (x"74",x"4b",x"49",x"6a"),
  1762 => (x"c2",x"9b",x"c3",x"2b"),
  1763 => (x"70",x"30",x"74",x"48"),
  1764 => (x"74",x"bc",x"ff",x"4c"),
  1765 => (x"70",x"98",x"71",x"48"),
  1766 => (x"87",x"d3",x"f6",x"7a"),
  1767 => (x"ef",x"fa",x"48",x"73"),
  1768 => (x"00",x"00",x"00",x"87"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"00",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"00",x"00"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"00",x"00",x"00",x"00"),
  1774 => (x"00",x"00",x"00",x"00"),
  1775 => (x"00",x"00",x"00",x"00"),
  1776 => (x"00",x"00",x"00",x"00"),
  1777 => (x"00",x"00",x"00",x"00"),
  1778 => (x"00",x"00",x"00",x"00"),
  1779 => (x"00",x"00",x"00",x"00"),
  1780 => (x"00",x"00",x"00",x"00"),
  1781 => (x"00",x"00",x"00",x"00"),
  1782 => (x"00",x"00",x"00",x"00"),
  1783 => (x"00",x"00",x"00",x"00"),
  1784 => (x"26",x"1e",x"16",x"00"),
  1785 => (x"3d",x"36",x"2e",x"25"),
  1786 => (x"d0",x"ff",x"1e",x"3e"),
  1787 => (x"78",x"e1",x"c8",x"48"),
  1788 => (x"d4",x"ff",x"48",x"71"),
  1789 => (x"66",x"c4",x"78",x"08"),
  1790 => (x"08",x"d4",x"ff",x"48"),
  1791 => (x"1e",x"4f",x"26",x"78"),
  1792 => (x"66",x"c4",x"4a",x"71"),
  1793 => (x"49",x"72",x"1e",x"49"),
  1794 => (x"ff",x"87",x"de",x"ff"),
  1795 => (x"e0",x"c0",x"48",x"d0"),
  1796 => (x"4f",x"26",x"26",x"78"),
  1797 => (x"c2",x"4a",x"71",x"1e"),
  1798 => (x"c3",x"03",x"aa",x"b7"),
  1799 => (x"87",x"c2",x"82",x"87"),
  1800 => (x"66",x"c4",x"82",x"ce"),
  1801 => (x"ff",x"49",x"72",x"1e"),
  1802 => (x"26",x"26",x"87",x"d5"),
  1803 => (x"d4",x"ff",x"1e",x"4f"),
  1804 => (x"7a",x"ff",x"c3",x"4a"),
  1805 => (x"c8",x"48",x"d0",x"ff"),
  1806 => (x"7a",x"de",x"78",x"e1"),
  1807 => (x"bf",x"dd",x"cc",x"c3"),
  1808 => (x"c8",x"48",x"49",x"7a"),
  1809 => (x"71",x"7a",x"70",x"28"),
  1810 => (x"70",x"28",x"d0",x"48"),
  1811 => (x"d8",x"48",x"71",x"7a"),
  1812 => (x"ff",x"7a",x"70",x"28"),
  1813 => (x"e0",x"c0",x"48",x"d0"),
  1814 => (x"0e",x"4f",x"26",x"78"),
  1815 => (x"5d",x"5c",x"5b",x"5e"),
  1816 => (x"c3",x"4c",x"71",x"0e"),
  1817 => (x"4d",x"bf",x"dd",x"cc"),
  1818 => (x"d0",x"2b",x"74",x"4b"),
  1819 => (x"83",x"c1",x"9b",x"66"),
  1820 => (x"04",x"ab",x"66",x"d4"),
  1821 => (x"4b",x"c0",x"87",x"c2"),
  1822 => (x"66",x"d0",x"4a",x"74"),
  1823 => (x"ff",x"31",x"72",x"49"),
  1824 => (x"73",x"99",x"75",x"b9"),
  1825 => (x"70",x"30",x"72",x"48"),
  1826 => (x"b0",x"71",x"48",x"4a"),
  1827 => (x"58",x"e1",x"cc",x"c3"),
  1828 => (x"26",x"87",x"da",x"fe"),
  1829 => (x"26",x"4c",x"26",x"4d"),
  1830 => (x"0e",x"4f",x"26",x"4b"),
  1831 => (x"5d",x"5c",x"5b",x"5e"),
  1832 => (x"4c",x"71",x"1e",x"0e"),
  1833 => (x"4b",x"e1",x"cc",x"c3"),
  1834 => (x"f4",x"c0",x"4a",x"c0"),
  1835 => (x"d4",x"d0",x"fe",x"49"),
  1836 => (x"c3",x"1e",x"74",x"87"),
  1837 => (x"fe",x"49",x"e1",x"cc"),
  1838 => (x"c4",x"87",x"cc",x"ee"),
  1839 => (x"02",x"98",x"70",x"86"),
  1840 => (x"c4",x"87",x"ea",x"c0"),
  1841 => (x"1e",x"4d",x"a6",x"1e"),
  1842 => (x"49",x"e1",x"cc",x"c3"),
  1843 => (x"87",x"fd",x"f3",x"fe"),
  1844 => (x"98",x"70",x"86",x"c8"),
  1845 => (x"75",x"87",x"d6",x"02"),
  1846 => (x"e3",x"f4",x"c1",x"4a"),
  1847 => (x"fe",x"4b",x"c4",x"49"),
  1848 => (x"70",x"87",x"c7",x"ce"),
  1849 => (x"87",x"ca",x"02",x"98"),
  1850 => (x"ed",x"c0",x"48",x"c0"),
  1851 => (x"c0",x"48",x"c0",x"87"),
  1852 => (x"f3",x"c0",x"87",x"e8"),
  1853 => (x"87",x"c4",x"c1",x"87"),
  1854 => (x"c8",x"02",x"98",x"70"),
  1855 => (x"87",x"fc",x"c0",x"87"),
  1856 => (x"f8",x"05",x"98",x"70"),
  1857 => (x"c1",x"cd",x"c3",x"87"),
  1858 => (x"87",x"cc",x"02",x"bf"),
  1859 => (x"48",x"dd",x"cc",x"c3"),
  1860 => (x"bf",x"c1",x"cd",x"c3"),
  1861 => (x"87",x"d5",x"fc",x"78"),
  1862 => (x"26",x"26",x"48",x"c1"),
  1863 => (x"26",x"4c",x"26",x"4d"),
  1864 => (x"5b",x"4f",x"26",x"4b"),
  1865 => (x"00",x"43",x"52",x"41"),
  1866 => (x"c3",x"1e",x"c0",x"1e"),
  1867 => (x"fe",x"49",x"e1",x"cc"),
  1868 => (x"c3",x"87",x"f3",x"f0"),
  1869 => (x"c0",x"48",x"f9",x"cc"),
  1870 => (x"4f",x"26",x"26",x"78"),
  1871 => (x"5c",x"5b",x"5e",x"0e"),
  1872 => (x"86",x"f4",x"0e",x"5d"),
  1873 => (x"c0",x"48",x"a6",x"c4"),
  1874 => (x"f9",x"cc",x"c3",x"78"),
  1875 => (x"b7",x"c3",x"48",x"bf"),
  1876 => (x"87",x"d1",x"03",x"a8"),
  1877 => (x"bf",x"f9",x"cc",x"c3"),
  1878 => (x"c3",x"80",x"c1",x"48"),
  1879 => (x"c0",x"58",x"fd",x"cc"),
  1880 => (x"e2",x"c6",x"48",x"fb"),
  1881 => (x"e1",x"cc",x"c3",x"87"),
  1882 => (x"f4",x"f5",x"fe",x"49"),
  1883 => (x"c3",x"4c",x"70",x"87"),
  1884 => (x"4a",x"bf",x"f9",x"cc"),
  1885 => (x"d8",x"02",x"8a",x"c3"),
  1886 => (x"02",x"8a",x"c1",x"87"),
  1887 => (x"8a",x"87",x"cb",x"c5"),
  1888 => (x"87",x"f6",x"c2",x"02"),
  1889 => (x"cd",x"c1",x"02",x"8a"),
  1890 => (x"c3",x"02",x"8a",x"87"),
  1891 => (x"e1",x"c5",x"87",x"e2"),
  1892 => (x"75",x"4d",x"c0",x"87"),
  1893 => (x"c1",x"92",x"c4",x"4a"),
  1894 => (x"c3",x"82",x"e5",x"fc"),
  1895 => (x"75",x"48",x"f5",x"cc"),
  1896 => (x"6e",x"7e",x"70",x"80"),
  1897 => (x"49",x"4b",x"bf",x"97"),
  1898 => (x"c1",x"48",x"6e",x"4b"),
  1899 => (x"81",x"6a",x"50",x"a3"),
  1900 => (x"a6",x"cc",x"48",x"11"),
  1901 => (x"02",x"ac",x"70",x"58"),
  1902 => (x"48",x"6e",x"87",x"c4"),
  1903 => (x"66",x"c8",x"50",x"c0"),
  1904 => (x"c3",x"87",x"c7",x"05"),
  1905 => (x"c4",x"48",x"f9",x"cc"),
  1906 => (x"85",x"c1",x"78",x"a5"),
  1907 => (x"04",x"ad",x"b7",x"c4"),
  1908 => (x"c4",x"87",x"c0",x"ff"),
  1909 => (x"cd",x"c3",x"87",x"dc"),
  1910 => (x"c8",x"48",x"bf",x"c5"),
  1911 => (x"d1",x"01",x"a8",x"b7"),
  1912 => (x"02",x"ac",x"ca",x"87"),
  1913 => (x"ac",x"cd",x"87",x"cc"),
  1914 => (x"c0",x"87",x"c7",x"02"),
  1915 => (x"c0",x"03",x"ac",x"b7"),
  1916 => (x"cd",x"c3",x"87",x"f3"),
  1917 => (x"c8",x"4b",x"bf",x"c5"),
  1918 => (x"d2",x"03",x"ab",x"b7"),
  1919 => (x"c9",x"cd",x"c3",x"87"),
  1920 => (x"c0",x"81",x"73",x"49"),
  1921 => (x"83",x"c1",x"51",x"e0"),
  1922 => (x"04",x"ab",x"b7",x"c8"),
  1923 => (x"c3",x"87",x"ee",x"ff"),
  1924 => (x"c1",x"48",x"d1",x"cd"),
  1925 => (x"cf",x"c1",x"50",x"d2"),
  1926 => (x"50",x"cd",x"c1",x"50"),
  1927 => (x"80",x"e4",x"50",x"c0"),
  1928 => (x"cd",x"c3",x"78",x"c3"),
  1929 => (x"c5",x"cd",x"c3",x"87"),
  1930 => (x"c1",x"48",x"49",x"bf"),
  1931 => (x"c9",x"cd",x"c3",x"80"),
  1932 => (x"a0",x"c4",x"48",x"58"),
  1933 => (x"c2",x"51",x"74",x"81"),
  1934 => (x"f0",x"c0",x"87",x"f8"),
  1935 => (x"da",x"04",x"ac",x"b7"),
  1936 => (x"b7",x"f9",x"c0",x"87"),
  1937 => (x"87",x"d3",x"01",x"ac"),
  1938 => (x"bf",x"fd",x"cc",x"c3"),
  1939 => (x"74",x"91",x"ca",x"49"),
  1940 => (x"8a",x"f0",x"c0",x"4a"),
  1941 => (x"48",x"fd",x"cc",x"c3"),
  1942 => (x"ca",x"78",x"a1",x"72"),
  1943 => (x"c6",x"c0",x"02",x"ac"),
  1944 => (x"05",x"ac",x"cd",x"87"),
  1945 => (x"c3",x"87",x"cb",x"c2"),
  1946 => (x"c3",x"48",x"f9",x"cc"),
  1947 => (x"87",x"c2",x"c2",x"78"),
  1948 => (x"ac",x"b7",x"f0",x"c0"),
  1949 => (x"c0",x"87",x"db",x"04"),
  1950 => (x"01",x"ac",x"b7",x"f9"),
  1951 => (x"c3",x"87",x"d3",x"c0"),
  1952 => (x"49",x"bf",x"c1",x"cd"),
  1953 => (x"4a",x"74",x"91",x"d0"),
  1954 => (x"c3",x"8a",x"f0",x"c0"),
  1955 => (x"72",x"48",x"c1",x"cd"),
  1956 => (x"c1",x"c1",x"78",x"a1"),
  1957 => (x"c0",x"04",x"ac",x"b7"),
  1958 => (x"c6",x"c1",x"87",x"db"),
  1959 => (x"c0",x"01",x"ac",x"b7"),
  1960 => (x"cd",x"c3",x"87",x"d3"),
  1961 => (x"d0",x"49",x"bf",x"c1"),
  1962 => (x"c0",x"4a",x"74",x"91"),
  1963 => (x"cd",x"c3",x"8a",x"f7"),
  1964 => (x"a1",x"72",x"48",x"c1"),
  1965 => (x"02",x"ac",x"ca",x"78"),
  1966 => (x"cd",x"87",x"c6",x"c0"),
  1967 => (x"f1",x"c0",x"05",x"ac"),
  1968 => (x"f9",x"cc",x"c3",x"87"),
  1969 => (x"c0",x"78",x"c3",x"48"),
  1970 => (x"e2",x"c0",x"87",x"e8"),
  1971 => (x"c9",x"c0",x"05",x"ac"),
  1972 => (x"48",x"a6",x"c4",x"87"),
  1973 => (x"c0",x"78",x"fb",x"c0"),
  1974 => (x"ac",x"ca",x"87",x"d8"),
  1975 => (x"87",x"c6",x"c0",x"02"),
  1976 => (x"c0",x"05",x"ac",x"cd"),
  1977 => (x"cc",x"c3",x"87",x"c9"),
  1978 => (x"78",x"c3",x"48",x"f9"),
  1979 => (x"c8",x"87",x"c3",x"c0"),
  1980 => (x"b7",x"c0",x"5c",x"a6"),
  1981 => (x"c4",x"c0",x"03",x"ac"),
  1982 => (x"ca",x"c0",x"48",x"87"),
  1983 => (x"02",x"66",x"c4",x"87"),
  1984 => (x"48",x"87",x"c6",x"f9"),
  1985 => (x"f4",x"99",x"ff",x"c3"),
  1986 => (x"87",x"cf",x"f8",x"8e"),
  1987 => (x"46",x"4e",x"4f",x"43"),
  1988 => (x"4f",x"4d",x"00",x"3d"),
  1989 => (x"41",x"4e",x"00",x"44"),
  1990 => (x"44",x"00",x"45",x"4d"),
  1991 => (x"55",x"41",x"46",x"45"),
  1992 => (x"30",x"3d",x"54",x"4c"),
  1993 => (x"00",x"1f",x"0c",x"00"),
  1994 => (x"00",x"1f",x"12",x"00"),
  1995 => (x"00",x"1f",x"16",x"00"),
  1996 => (x"00",x"1f",x"1b",x"00"),
  1997 => (x"d0",x"ff",x"1e",x"00"),
  1998 => (x"78",x"c9",x"c8",x"48"),
  1999 => (x"d4",x"ff",x"48",x"71"),
  2000 => (x"4f",x"26",x"78",x"08"),
  2001 => (x"49",x"4a",x"71",x"1e"),
  2002 => (x"d0",x"ff",x"87",x"eb"),
  2003 => (x"26",x"78",x"c8",x"48"),
  2004 => (x"1e",x"73",x"1e",x"4f"),
  2005 => (x"cd",x"c3",x"4b",x"71"),
  2006 => (x"c3",x"02",x"bf",x"e1"),
  2007 => (x"87",x"eb",x"c2",x"87"),
  2008 => (x"c8",x"48",x"d0",x"ff"),
  2009 => (x"49",x"73",x"78",x"c9"),
  2010 => (x"ff",x"b1",x"e0",x"c0"),
  2011 => (x"78",x"71",x"48",x"d4"),
  2012 => (x"48",x"d5",x"cd",x"c3"),
  2013 => (x"66",x"c8",x"78",x"c0"),
  2014 => (x"c3",x"87",x"c5",x"02"),
  2015 => (x"87",x"c2",x"49",x"ff"),
  2016 => (x"cd",x"c3",x"49",x"c0"),
  2017 => (x"66",x"cc",x"59",x"dd"),
  2018 => (x"c5",x"87",x"c6",x"02"),
  2019 => (x"c4",x"4a",x"d5",x"d5"),
  2020 => (x"ff",x"ff",x"cf",x"87"),
  2021 => (x"e1",x"cd",x"c3",x"4a"),
  2022 => (x"e1",x"cd",x"c3",x"5a"),
  2023 => (x"c4",x"78",x"c1",x"48"),
  2024 => (x"26",x"4d",x"26",x"87"),
  2025 => (x"26",x"4b",x"26",x"4c"),
  2026 => (x"5b",x"5e",x"0e",x"4f"),
  2027 => (x"71",x"0e",x"5d",x"5c"),
  2028 => (x"dd",x"cd",x"c3",x"4a"),
  2029 => (x"9a",x"72",x"4c",x"bf"),
  2030 => (x"49",x"87",x"cb",x"02"),
  2031 => (x"fd",x"c1",x"91",x"c8"),
  2032 => (x"83",x"71",x"4b",x"c7"),
  2033 => (x"c1",x"c2",x"87",x"c4"),
  2034 => (x"4d",x"c0",x"4b",x"c7"),
  2035 => (x"99",x"74",x"49",x"13"),
  2036 => (x"bf",x"d9",x"cd",x"c3"),
  2037 => (x"48",x"d4",x"ff",x"b9"),
  2038 => (x"b7",x"c1",x"78",x"71"),
  2039 => (x"b7",x"c8",x"85",x"2c"),
  2040 => (x"87",x"e8",x"04",x"ad"),
  2041 => (x"bf",x"d5",x"cd",x"c3"),
  2042 => (x"c3",x"80",x"c8",x"48"),
  2043 => (x"fe",x"58",x"d9",x"cd"),
  2044 => (x"73",x"1e",x"87",x"ef"),
  2045 => (x"13",x"4b",x"71",x"1e"),
  2046 => (x"cb",x"02",x"9a",x"4a"),
  2047 => (x"fe",x"49",x"72",x"87"),
  2048 => (x"4a",x"13",x"87",x"e7"),
  2049 => (x"87",x"f5",x"05",x"9a"),
  2050 => (x"1e",x"87",x"da",x"fe"),
  2051 => (x"bf",x"d5",x"cd",x"c3"),
  2052 => (x"d5",x"cd",x"c3",x"49"),
  2053 => (x"78",x"a1",x"c1",x"48"),
  2054 => (x"a9",x"b7",x"c0",x"c4"),
  2055 => (x"ff",x"87",x"db",x"03"),
  2056 => (x"cd",x"c3",x"48",x"d4"),
  2057 => (x"c3",x"78",x"bf",x"d9"),
  2058 => (x"49",x"bf",x"d5",x"cd"),
  2059 => (x"48",x"d5",x"cd",x"c3"),
  2060 => (x"c4",x"78",x"a1",x"c1"),
  2061 => (x"04",x"a9",x"b7",x"c0"),
  2062 => (x"d0",x"ff",x"87",x"e5"),
  2063 => (x"c3",x"78",x"c8",x"48"),
  2064 => (x"c0",x"48",x"e1",x"cd"),
  2065 => (x"00",x"4f",x"26",x"78"),
  2066 => (x"00",x"00",x"00",x"00"),
  2067 => (x"00",x"00",x"00",x"00"),
  2068 => (x"5f",x"5f",x"00",x"00"),
  2069 => (x"00",x"00",x"00",x"00"),
  2070 => (x"03",x"00",x"03",x"03"),
  2071 => (x"14",x"00",x"00",x"03"),
  2072 => (x"7f",x"14",x"7f",x"7f"),
  2073 => (x"00",x"00",x"14",x"7f"),
  2074 => (x"6b",x"6b",x"2e",x"24"),
  2075 => (x"4c",x"00",x"12",x"3a"),
  2076 => (x"6c",x"18",x"36",x"6a"),
  2077 => (x"30",x"00",x"32",x"56"),
  2078 => (x"77",x"59",x"4f",x"7e"),
  2079 => (x"00",x"40",x"68",x"3a"),
  2080 => (x"03",x"07",x"04",x"00"),
  2081 => (x"00",x"00",x"00",x"00"),
  2082 => (x"63",x"3e",x"1c",x"00"),
  2083 => (x"00",x"00",x"00",x"41"),
  2084 => (x"3e",x"63",x"41",x"00"),
  2085 => (x"08",x"00",x"00",x"1c"),
  2086 => (x"1c",x"1c",x"3e",x"2a"),
  2087 => (x"00",x"08",x"2a",x"3e"),
  2088 => (x"3e",x"3e",x"08",x"08"),
  2089 => (x"00",x"00",x"08",x"08"),
  2090 => (x"60",x"e0",x"80",x"00"),
  2091 => (x"00",x"00",x"00",x"00"),
  2092 => (x"08",x"08",x"08",x"08"),
  2093 => (x"00",x"00",x"08",x"08"),
  2094 => (x"60",x"60",x"00",x"00"),
  2095 => (x"40",x"00",x"00",x"00"),
  2096 => (x"0c",x"18",x"30",x"60"),
  2097 => (x"00",x"01",x"03",x"06"),
  2098 => (x"4d",x"59",x"7f",x"3e"),
  2099 => (x"00",x"00",x"3e",x"7f"),
  2100 => (x"7f",x"7f",x"06",x"04"),
  2101 => (x"00",x"00",x"00",x"00"),
  2102 => (x"59",x"71",x"63",x"42"),
  2103 => (x"00",x"00",x"46",x"4f"),
  2104 => (x"49",x"49",x"63",x"22"),
  2105 => (x"18",x"00",x"36",x"7f"),
  2106 => (x"7f",x"13",x"16",x"1c"),
  2107 => (x"00",x"00",x"10",x"7f"),
  2108 => (x"45",x"45",x"67",x"27"),
  2109 => (x"00",x"00",x"39",x"7d"),
  2110 => (x"49",x"4b",x"7e",x"3c"),
  2111 => (x"00",x"00",x"30",x"79"),
  2112 => (x"79",x"71",x"01",x"01"),
  2113 => (x"00",x"00",x"07",x"0f"),
  2114 => (x"49",x"49",x"7f",x"36"),
  2115 => (x"00",x"00",x"36",x"7f"),
  2116 => (x"69",x"49",x"4f",x"06"),
  2117 => (x"00",x"00",x"1e",x"3f"),
  2118 => (x"66",x"66",x"00",x"00"),
  2119 => (x"00",x"00",x"00",x"00"),
  2120 => (x"66",x"e6",x"80",x"00"),
  2121 => (x"00",x"00",x"00",x"00"),
  2122 => (x"14",x"14",x"08",x"08"),
  2123 => (x"00",x"00",x"22",x"22"),
  2124 => (x"14",x"14",x"14",x"14"),
  2125 => (x"00",x"00",x"14",x"14"),
  2126 => (x"14",x"14",x"22",x"22"),
  2127 => (x"00",x"00",x"08",x"08"),
  2128 => (x"59",x"51",x"03",x"02"),
  2129 => (x"3e",x"00",x"06",x"0f"),
  2130 => (x"55",x"5d",x"41",x"7f"),
  2131 => (x"00",x"00",x"1e",x"1f"),
  2132 => (x"09",x"09",x"7f",x"7e"),
  2133 => (x"00",x"00",x"7e",x"7f"),
  2134 => (x"49",x"49",x"7f",x"7f"),
  2135 => (x"00",x"00",x"36",x"7f"),
  2136 => (x"41",x"63",x"3e",x"1c"),
  2137 => (x"00",x"00",x"41",x"41"),
  2138 => (x"63",x"41",x"7f",x"7f"),
  2139 => (x"00",x"00",x"1c",x"3e"),
  2140 => (x"49",x"49",x"7f",x"7f"),
  2141 => (x"00",x"00",x"41",x"41"),
  2142 => (x"09",x"09",x"7f",x"7f"),
  2143 => (x"00",x"00",x"01",x"01"),
  2144 => (x"49",x"41",x"7f",x"3e"),
  2145 => (x"00",x"00",x"7a",x"7b"),
  2146 => (x"08",x"08",x"7f",x"7f"),
  2147 => (x"00",x"00",x"7f",x"7f"),
  2148 => (x"7f",x"7f",x"41",x"00"),
  2149 => (x"00",x"00",x"00",x"41"),
  2150 => (x"40",x"40",x"60",x"20"),
  2151 => (x"7f",x"00",x"3f",x"7f"),
  2152 => (x"36",x"1c",x"08",x"7f"),
  2153 => (x"00",x"00",x"41",x"63"),
  2154 => (x"40",x"40",x"7f",x"7f"),
  2155 => (x"7f",x"00",x"40",x"40"),
  2156 => (x"06",x"0c",x"06",x"7f"),
  2157 => (x"7f",x"00",x"7f",x"7f"),
  2158 => (x"18",x"0c",x"06",x"7f"),
  2159 => (x"00",x"00",x"7f",x"7f"),
  2160 => (x"41",x"41",x"7f",x"3e"),
  2161 => (x"00",x"00",x"3e",x"7f"),
  2162 => (x"09",x"09",x"7f",x"7f"),
  2163 => (x"3e",x"00",x"06",x"0f"),
  2164 => (x"7f",x"61",x"41",x"7f"),
  2165 => (x"00",x"00",x"40",x"7e"),
  2166 => (x"19",x"09",x"7f",x"7f"),
  2167 => (x"00",x"00",x"66",x"7f"),
  2168 => (x"59",x"4d",x"6f",x"26"),
  2169 => (x"00",x"00",x"32",x"7b"),
  2170 => (x"7f",x"7f",x"01",x"01"),
  2171 => (x"00",x"00",x"01",x"01"),
  2172 => (x"40",x"40",x"7f",x"3f"),
  2173 => (x"00",x"00",x"3f",x"7f"),
  2174 => (x"70",x"70",x"3f",x"0f"),
  2175 => (x"7f",x"00",x"0f",x"3f"),
  2176 => (x"30",x"18",x"30",x"7f"),
  2177 => (x"41",x"00",x"7f",x"7f"),
  2178 => (x"1c",x"1c",x"36",x"63"),
  2179 => (x"01",x"41",x"63",x"36"),
  2180 => (x"7c",x"7c",x"06",x"03"),
  2181 => (x"61",x"01",x"03",x"06"),
  2182 => (x"47",x"4d",x"59",x"71"),
  2183 => (x"00",x"00",x"41",x"43"),
  2184 => (x"41",x"7f",x"7f",x"00"),
  2185 => (x"01",x"00",x"00",x"41"),
  2186 => (x"18",x"0c",x"06",x"03"),
  2187 => (x"00",x"40",x"60",x"30"),
  2188 => (x"7f",x"41",x"41",x"00"),
  2189 => (x"08",x"00",x"00",x"7f"),
  2190 => (x"06",x"03",x"06",x"0c"),
  2191 => (x"80",x"00",x"08",x"0c"),
  2192 => (x"80",x"80",x"80",x"80"),
  2193 => (x"00",x"00",x"80",x"80"),
  2194 => (x"07",x"03",x"00",x"00"),
  2195 => (x"00",x"00",x"00",x"04"),
  2196 => (x"54",x"54",x"74",x"20"),
  2197 => (x"00",x"00",x"78",x"7c"),
  2198 => (x"44",x"44",x"7f",x"7f"),
  2199 => (x"00",x"00",x"38",x"7c"),
  2200 => (x"44",x"44",x"7c",x"38"),
  2201 => (x"00",x"00",x"00",x"44"),
  2202 => (x"44",x"44",x"7c",x"38"),
  2203 => (x"00",x"00",x"7f",x"7f"),
  2204 => (x"54",x"54",x"7c",x"38"),
  2205 => (x"00",x"00",x"18",x"5c"),
  2206 => (x"05",x"7f",x"7e",x"04"),
  2207 => (x"00",x"00",x"00",x"05"),
  2208 => (x"a4",x"a4",x"bc",x"18"),
  2209 => (x"00",x"00",x"7c",x"fc"),
  2210 => (x"04",x"04",x"7f",x"7f"),
  2211 => (x"00",x"00",x"78",x"7c"),
  2212 => (x"7d",x"3d",x"00",x"00"),
  2213 => (x"00",x"00",x"00",x"40"),
  2214 => (x"fd",x"80",x"80",x"80"),
  2215 => (x"00",x"00",x"00",x"7d"),
  2216 => (x"38",x"10",x"7f",x"7f"),
  2217 => (x"00",x"00",x"44",x"6c"),
  2218 => (x"7f",x"3f",x"00",x"00"),
  2219 => (x"7c",x"00",x"00",x"40"),
  2220 => (x"0c",x"18",x"0c",x"7c"),
  2221 => (x"00",x"00",x"78",x"7c"),
  2222 => (x"04",x"04",x"7c",x"7c"),
  2223 => (x"00",x"00",x"78",x"7c"),
  2224 => (x"44",x"44",x"7c",x"38"),
  2225 => (x"00",x"00",x"38",x"7c"),
  2226 => (x"24",x"24",x"fc",x"fc"),
  2227 => (x"00",x"00",x"18",x"3c"),
  2228 => (x"24",x"24",x"3c",x"18"),
  2229 => (x"00",x"00",x"fc",x"fc"),
  2230 => (x"04",x"04",x"7c",x"7c"),
  2231 => (x"00",x"00",x"08",x"0c"),
  2232 => (x"54",x"54",x"5c",x"48"),
  2233 => (x"00",x"00",x"20",x"74"),
  2234 => (x"44",x"7f",x"3f",x"04"),
  2235 => (x"00",x"00",x"00",x"44"),
  2236 => (x"40",x"40",x"7c",x"3c"),
  2237 => (x"00",x"00",x"7c",x"7c"),
  2238 => (x"60",x"60",x"3c",x"1c"),
  2239 => (x"3c",x"00",x"1c",x"3c"),
  2240 => (x"60",x"30",x"60",x"7c"),
  2241 => (x"44",x"00",x"3c",x"7c"),
  2242 => (x"38",x"10",x"38",x"6c"),
  2243 => (x"00",x"00",x"44",x"6c"),
  2244 => (x"60",x"e0",x"bc",x"1c"),
  2245 => (x"00",x"00",x"1c",x"3c"),
  2246 => (x"5c",x"74",x"64",x"44"),
  2247 => (x"00",x"00",x"44",x"4c"),
  2248 => (x"77",x"3e",x"08",x"08"),
  2249 => (x"00",x"00",x"41",x"41"),
  2250 => (x"7f",x"7f",x"00",x"00"),
  2251 => (x"00",x"00",x"00",x"00"),
  2252 => (x"3e",x"77",x"41",x"41"),
  2253 => (x"02",x"00",x"08",x"08"),
  2254 => (x"02",x"03",x"01",x"01"),
  2255 => (x"7f",x"00",x"01",x"02"),
  2256 => (x"7f",x"7f",x"7f",x"7f"),
  2257 => (x"08",x"00",x"7f",x"7f"),
  2258 => (x"3e",x"1c",x"1c",x"08"),
  2259 => (x"7f",x"7f",x"7f",x"3e"),
  2260 => (x"1c",x"3e",x"3e",x"7f"),
  2261 => (x"00",x"08",x"08",x"1c"),
  2262 => (x"7c",x"7c",x"18",x"10"),
  2263 => (x"00",x"00",x"10",x"18"),
  2264 => (x"7c",x"7c",x"30",x"10"),
  2265 => (x"10",x"00",x"10",x"30"),
  2266 => (x"78",x"60",x"60",x"30"),
  2267 => (x"42",x"00",x"06",x"1e"),
  2268 => (x"3c",x"18",x"3c",x"66"),
  2269 => (x"78",x"00",x"42",x"66"),
  2270 => (x"c6",x"c2",x"6a",x"38"),
  2271 => (x"60",x"00",x"38",x"6c"),
  2272 => (x"00",x"60",x"00",x"00"),
  2273 => (x"0e",x"00",x"60",x"00"),
  2274 => (x"5d",x"5c",x"5b",x"5e"),
  2275 => (x"4c",x"71",x"1e",x"0e"),
  2276 => (x"bf",x"f2",x"cd",x"c3"),
  2277 => (x"c0",x"4b",x"c0",x"4d"),
  2278 => (x"02",x"ab",x"74",x"1e"),
  2279 => (x"a6",x"c4",x"87",x"c7"),
  2280 => (x"c5",x"78",x"c0",x"48"),
  2281 => (x"48",x"a6",x"c4",x"87"),
  2282 => (x"66",x"c4",x"78",x"c1"),
  2283 => (x"ee",x"49",x"73",x"1e"),
  2284 => (x"86",x"c8",x"87",x"df"),
  2285 => (x"ef",x"49",x"e0",x"c0"),
  2286 => (x"a5",x"c4",x"87",x"ef"),
  2287 => (x"f0",x"49",x"6a",x"4a"),
  2288 => (x"c6",x"f1",x"87",x"f0"),
  2289 => (x"c1",x"85",x"cb",x"87"),
  2290 => (x"ab",x"b7",x"c8",x"83"),
  2291 => (x"87",x"c7",x"ff",x"04"),
  2292 => (x"26",x"4d",x"26",x"26"),
  2293 => (x"26",x"4b",x"26",x"4c"),
  2294 => (x"4a",x"71",x"1e",x"4f"),
  2295 => (x"5a",x"f6",x"cd",x"c3"),
  2296 => (x"48",x"f6",x"cd",x"c3"),
  2297 => (x"fe",x"49",x"78",x"c7"),
  2298 => (x"4f",x"26",x"87",x"dd"),
  2299 => (x"71",x"1e",x"73",x"1e"),
  2300 => (x"aa",x"b7",x"c0",x"4a"),
  2301 => (x"c2",x"87",x"d3",x"03"),
  2302 => (x"05",x"bf",x"c2",x"e0"),
  2303 => (x"4b",x"c1",x"87",x"c4"),
  2304 => (x"4b",x"c0",x"87",x"c2"),
  2305 => (x"5b",x"c6",x"e0",x"c2"),
  2306 => (x"e0",x"c2",x"87",x"c4"),
  2307 => (x"e0",x"c2",x"5a",x"c6"),
  2308 => (x"c1",x"4a",x"bf",x"c2"),
  2309 => (x"a2",x"c0",x"c1",x"9a"),
  2310 => (x"87",x"e8",x"ec",x"49"),
  2311 => (x"bf",x"ea",x"df",x"c2"),
  2312 => (x"c2",x"e0",x"c2",x"49"),
  2313 => (x"48",x"fc",x"b1",x"bf"),
  2314 => (x"e8",x"fe",x"78",x"71"),
  2315 => (x"4a",x"71",x"1e",x"87"),
  2316 => (x"72",x"1e",x"66",x"c4"),
  2317 => (x"db",x"df",x"ff",x"49"),
  2318 => (x"4f",x"26",x"26",x"87"),
  2319 => (x"c2",x"e0",x"c2",x"1e"),
  2320 => (x"e2",x"c0",x"49",x"bf"),
  2321 => (x"cd",x"c3",x"87",x"f0"),
  2322 => (x"bf",x"e8",x"48",x"ea"),
  2323 => (x"e6",x"cd",x"c3",x"78"),
  2324 => (x"78",x"bf",x"ec",x"48"),
  2325 => (x"bf",x"ea",x"cd",x"c3"),
  2326 => (x"ff",x"c3",x"49",x"4a"),
  2327 => (x"2a",x"b7",x"c8",x"99"),
  2328 => (x"b0",x"71",x"48",x"72"),
  2329 => (x"58",x"f2",x"cd",x"c3"),
  2330 => (x"5e",x"0e",x"4f",x"26"),
  2331 => (x"0e",x"5d",x"5c",x"5b"),
  2332 => (x"c7",x"ff",x"4b",x"71"),
  2333 => (x"e5",x"cd",x"c3",x"87"),
  2334 => (x"73",x"50",x"c0",x"48"),
  2335 => (x"e8",x"db",x"ff",x"49"),
  2336 => (x"4c",x"49",x"70",x"87"),
  2337 => (x"ee",x"cb",x"9c",x"c2"),
  2338 => (x"87",x"fe",x"cd",x"49"),
  2339 => (x"c3",x"4d",x"49",x"70"),
  2340 => (x"bf",x"97",x"e5",x"cd"),
  2341 => (x"87",x"e4",x"c1",x"05"),
  2342 => (x"c3",x"49",x"66",x"d0"),
  2343 => (x"99",x"bf",x"ee",x"cd"),
  2344 => (x"d4",x"87",x"d7",x"05"),
  2345 => (x"cd",x"c3",x"49",x"66"),
  2346 => (x"05",x"99",x"bf",x"e6"),
  2347 => (x"49",x"73",x"87",x"cc"),
  2348 => (x"87",x"f5",x"da",x"ff"),
  2349 => (x"c1",x"02",x"98",x"70"),
  2350 => (x"4c",x"c1",x"87",x"c2"),
  2351 => (x"75",x"87",x"fd",x"fd"),
  2352 => (x"87",x"d2",x"cd",x"49"),
  2353 => (x"c6",x"02",x"98",x"70"),
  2354 => (x"e5",x"cd",x"c3",x"87"),
  2355 => (x"c3",x"50",x"c1",x"48"),
  2356 => (x"bf",x"97",x"e5",x"cd"),
  2357 => (x"87",x"e4",x"c0",x"05"),
  2358 => (x"bf",x"ee",x"cd",x"c3"),
  2359 => (x"99",x"66",x"d0",x"49"),
  2360 => (x"87",x"d6",x"ff",x"05"),
  2361 => (x"bf",x"e6",x"cd",x"c3"),
  2362 => (x"99",x"66",x"d4",x"49"),
  2363 => (x"87",x"ca",x"ff",x"05"),
  2364 => (x"d9",x"ff",x"49",x"73"),
  2365 => (x"98",x"70",x"87",x"f3"),
  2366 => (x"87",x"fe",x"fe",x"05"),
  2367 => (x"d0",x"fb",x"48",x"74"),
  2368 => (x"5b",x"5e",x"0e",x"87"),
  2369 => (x"f8",x"0e",x"5d",x"5c"),
  2370 => (x"4c",x"4d",x"c0",x"86"),
  2371 => (x"c4",x"7e",x"bf",x"ec"),
  2372 => (x"cd",x"c3",x"48",x"a6"),
  2373 => (x"c0",x"78",x"bf",x"f2"),
  2374 => (x"f7",x"c1",x"1e",x"1e"),
  2375 => (x"87",x"ca",x"fd",x"49"),
  2376 => (x"98",x"70",x"86",x"c8"),
  2377 => (x"87",x"f3",x"c0",x"02"),
  2378 => (x"bf",x"ea",x"df",x"c2"),
  2379 => (x"c1",x"87",x"c4",x"05"),
  2380 => (x"c0",x"87",x"c2",x"7e"),
  2381 => (x"ea",x"df",x"c2",x"7e"),
  2382 => (x"ca",x"78",x"6e",x"48"),
  2383 => (x"66",x"c4",x"1e",x"fc"),
  2384 => (x"c4",x"87",x"c9",x"02"),
  2385 => (x"de",x"c2",x"48",x"a6"),
  2386 => (x"87",x"c7",x"78",x"c1"),
  2387 => (x"c2",x"48",x"a6",x"c4"),
  2388 => (x"c4",x"78",x"cc",x"de"),
  2389 => (x"ff",x"c8",x"49",x"66"),
  2390 => (x"c1",x"86",x"c4",x"87"),
  2391 => (x"c7",x"1e",x"c0",x"1e"),
  2392 => (x"87",x"c6",x"fc",x"49"),
  2393 => (x"98",x"70",x"86",x"c8"),
  2394 => (x"ff",x"87",x"ce",x"02"),
  2395 => (x"87",x"fc",x"f9",x"49"),
  2396 => (x"ff",x"49",x"da",x"c1"),
  2397 => (x"c1",x"87",x"f2",x"d7"),
  2398 => (x"e5",x"cd",x"c3",x"4d"),
  2399 => (x"c3",x"02",x"bf",x"97"),
  2400 => (x"87",x"e4",x"cf",x"87"),
  2401 => (x"bf",x"ea",x"cd",x"c3"),
  2402 => (x"c2",x"e0",x"c2",x"4b"),
  2403 => (x"e4",x"c1",x"05",x"bf"),
  2404 => (x"ea",x"df",x"c2",x"87"),
  2405 => (x"f1",x"c0",x"02",x"bf"),
  2406 => (x"48",x"a6",x"c4",x"87"),
  2407 => (x"78",x"c0",x"c0",x"c8"),
  2408 => (x"7e",x"ee",x"df",x"c2"),
  2409 => (x"49",x"bf",x"97",x"6e"),
  2410 => (x"80",x"c1",x"48",x"6e"),
  2411 => (x"ff",x"71",x"7e",x"70"),
  2412 => (x"70",x"87",x"f6",x"d6"),
  2413 => (x"87",x"c3",x"02",x"98"),
  2414 => (x"c4",x"b3",x"66",x"c4"),
  2415 => (x"b7",x"c1",x"48",x"66"),
  2416 => (x"58",x"a6",x"c8",x"28"),
  2417 => (x"ff",x"05",x"98",x"70"),
  2418 => (x"fd",x"c3",x"87",x"da"),
  2419 => (x"d8",x"d6",x"ff",x"49"),
  2420 => (x"49",x"fa",x"c3",x"87"),
  2421 => (x"87",x"d1",x"d6",x"ff"),
  2422 => (x"ff",x"c3",x"49",x"73"),
  2423 => (x"c0",x"1e",x"71",x"99"),
  2424 => (x"87",x"c9",x"f9",x"49"),
  2425 => (x"b7",x"c8",x"49",x"73"),
  2426 => (x"c1",x"1e",x"71",x"29"),
  2427 => (x"87",x"fd",x"f8",x"49"),
  2428 => (x"c7",x"c6",x"86",x"c8"),
  2429 => (x"ee",x"cd",x"c3",x"87"),
  2430 => (x"02",x"9b",x"4b",x"bf"),
  2431 => (x"df",x"c2",x"87",x"df"),
  2432 => (x"c8",x"49",x"bf",x"fe"),
  2433 => (x"98",x"70",x"87",x"d0"),
  2434 => (x"87",x"c4",x"c0",x"05"),
  2435 => (x"87",x"d3",x"4b",x"c0"),
  2436 => (x"c7",x"49",x"e0",x"c2"),
  2437 => (x"e0",x"c2",x"87",x"f4"),
  2438 => (x"c6",x"c0",x"58",x"c2"),
  2439 => (x"fe",x"df",x"c2",x"87"),
  2440 => (x"73",x"78",x"c0",x"48"),
  2441 => (x"05",x"99",x"c2",x"49"),
  2442 => (x"c3",x"87",x"cf",x"c0"),
  2443 => (x"d4",x"ff",x"49",x"eb"),
  2444 => (x"49",x"70",x"87",x"f7"),
  2445 => (x"c0",x"02",x"99",x"c2"),
  2446 => (x"4c",x"fb",x"87",x"c2"),
  2447 => (x"99",x"c1",x"49",x"73"),
  2448 => (x"87",x"cf",x"c0",x"05"),
  2449 => (x"ff",x"49",x"f4",x"c3"),
  2450 => (x"70",x"87",x"de",x"d4"),
  2451 => (x"02",x"99",x"c2",x"49"),
  2452 => (x"fa",x"87",x"c2",x"c0"),
  2453 => (x"c8",x"49",x"73",x"4c"),
  2454 => (x"cf",x"c0",x"05",x"99"),
  2455 => (x"49",x"f5",x"c3",x"87"),
  2456 => (x"87",x"c5",x"d4",x"ff"),
  2457 => (x"99",x"c2",x"49",x"70"),
  2458 => (x"87",x"d6",x"c0",x"02"),
  2459 => (x"bf",x"f6",x"cd",x"c3"),
  2460 => (x"87",x"ca",x"c0",x"02"),
  2461 => (x"c3",x"88",x"c1",x"48"),
  2462 => (x"c0",x"58",x"fa",x"cd"),
  2463 => (x"4c",x"ff",x"87",x"c2"),
  2464 => (x"49",x"73",x"4d",x"c1"),
  2465 => (x"c0",x"05",x"99",x"c4"),
  2466 => (x"f2",x"c3",x"87",x"cf"),
  2467 => (x"d8",x"d3",x"ff",x"49"),
  2468 => (x"c2",x"49",x"70",x"87"),
  2469 => (x"dc",x"c0",x"02",x"99"),
  2470 => (x"f6",x"cd",x"c3",x"87"),
  2471 => (x"c7",x"48",x"7e",x"bf"),
  2472 => (x"c0",x"03",x"a8",x"b7"),
  2473 => (x"48",x"6e",x"87",x"cb"),
  2474 => (x"cd",x"c3",x"80",x"c1"),
  2475 => (x"c2",x"c0",x"58",x"fa"),
  2476 => (x"c1",x"4c",x"fe",x"87"),
  2477 => (x"49",x"fd",x"c3",x"4d"),
  2478 => (x"87",x"ed",x"d2",x"ff"),
  2479 => (x"99",x"c2",x"49",x"70"),
  2480 => (x"87",x"d5",x"c0",x"02"),
  2481 => (x"bf",x"f6",x"cd",x"c3"),
  2482 => (x"87",x"c9",x"c0",x"02"),
  2483 => (x"48",x"f6",x"cd",x"c3"),
  2484 => (x"c2",x"c0",x"78",x"c0"),
  2485 => (x"c1",x"4c",x"fd",x"87"),
  2486 => (x"49",x"fa",x"c3",x"4d"),
  2487 => (x"87",x"c9",x"d2",x"ff"),
  2488 => (x"99",x"c2",x"49",x"70"),
  2489 => (x"87",x"d9",x"c0",x"02"),
  2490 => (x"bf",x"f6",x"cd",x"c3"),
  2491 => (x"a8",x"b7",x"c7",x"48"),
  2492 => (x"87",x"c9",x"c0",x"03"),
  2493 => (x"48",x"f6",x"cd",x"c3"),
  2494 => (x"c2",x"c0",x"78",x"c7"),
  2495 => (x"c1",x"4c",x"fc",x"87"),
  2496 => (x"ac",x"b7",x"c0",x"4d"),
  2497 => (x"87",x"d5",x"c0",x"03"),
  2498 => (x"c1",x"48",x"66",x"c4"),
  2499 => (x"7e",x"70",x"80",x"d8"),
  2500 => (x"c0",x"02",x"bf",x"6e"),
  2501 => (x"bf",x"6e",x"87",x"c7"),
  2502 => (x"73",x"49",x"74",x"4b"),
  2503 => (x"c3",x"1e",x"c0",x"0f"),
  2504 => (x"da",x"c1",x"1e",x"f0"),
  2505 => (x"87",x"c2",x"f5",x"49"),
  2506 => (x"98",x"70",x"86",x"c8"),
  2507 => (x"87",x"d9",x"c0",x"02"),
  2508 => (x"bf",x"f6",x"cd",x"c3"),
  2509 => (x"cb",x"49",x"6e",x"7e"),
  2510 => (x"4a",x"66",x"c4",x"91"),
  2511 => (x"02",x"6a",x"82",x"71"),
  2512 => (x"6a",x"87",x"c6",x"c0"),
  2513 => (x"73",x"49",x"6e",x"4b"),
  2514 => (x"02",x"9d",x"75",x"0f"),
  2515 => (x"c3",x"87",x"c8",x"c0"),
  2516 => (x"49",x"bf",x"f6",x"cd"),
  2517 => (x"c2",x"87",x"f0",x"f0"),
  2518 => (x"02",x"bf",x"c6",x"e0"),
  2519 => (x"49",x"87",x"dd",x"c0"),
  2520 => (x"70",x"87",x"f3",x"c2"),
  2521 => (x"d3",x"c0",x"02",x"98"),
  2522 => (x"f6",x"cd",x"c3",x"87"),
  2523 => (x"d6",x"f0",x"49",x"bf"),
  2524 => (x"f1",x"49",x"c0",x"87"),
  2525 => (x"e0",x"c2",x"87",x"f6"),
  2526 => (x"78",x"c0",x"48",x"c6"),
  2527 => (x"d0",x"f1",x"8e",x"f8"),
  2528 => (x"79",x"6f",x"4a",x"87"),
  2529 => (x"73",x"79",x"65",x"6b"),
  2530 => (x"00",x"6e",x"6f",x"20"),
  2531 => (x"6b",x"79",x"6f",x"4a"),
  2532 => (x"20",x"73",x"79",x"65"),
  2533 => (x"00",x"66",x"66",x"6f"),
  2534 => (x"5c",x"5b",x"5e",x"0e"),
  2535 => (x"71",x"1e",x"0e",x"5d"),
  2536 => (x"f2",x"cd",x"c3",x"4c"),
  2537 => (x"cd",x"c1",x"49",x"bf"),
  2538 => (x"d1",x"c1",x"4d",x"a1"),
  2539 => (x"74",x"7e",x"69",x"81"),
  2540 => (x"87",x"cf",x"02",x"9c"),
  2541 => (x"74",x"4b",x"a5",x"c4"),
  2542 => (x"f2",x"cd",x"c3",x"7b"),
  2543 => (x"d8",x"f0",x"49",x"bf"),
  2544 => (x"74",x"7b",x"6e",x"87"),
  2545 => (x"87",x"c4",x"05",x"9c"),
  2546 => (x"87",x"c2",x"4b",x"c0"),
  2547 => (x"49",x"73",x"4b",x"c1"),
  2548 => (x"d4",x"87",x"d9",x"f0"),
  2549 => (x"87",x"c8",x"02",x"66"),
  2550 => (x"87",x"ee",x"c0",x"49"),
  2551 => (x"87",x"c2",x"4a",x"70"),
  2552 => (x"e0",x"c2",x"4a",x"c0"),
  2553 => (x"ef",x"26",x"5a",x"ca"),
  2554 => (x"00",x"00",x"87",x"e7"),
  2555 => (x"12",x"58",x"00",x"00"),
  2556 => (x"1b",x"1d",x"14",x"11"),
  2557 => (x"59",x"5a",x"23",x"1c"),
  2558 => (x"f2",x"f5",x"94",x"91"),
  2559 => (x"00",x"00",x"f4",x"eb"),
  2560 => (x"00",x"00",x"00",x"00"),
  2561 => (x"00",x"00",x"00",x"00"),
  2562 => (x"71",x"1e",x"00",x"00"),
  2563 => (x"bf",x"c8",x"ff",x"4a"),
  2564 => (x"48",x"a1",x"72",x"49"),
  2565 => (x"ff",x"1e",x"4f",x"26"),
  2566 => (x"fe",x"89",x"bf",x"c8"),
  2567 => (x"c0",x"c0",x"c0",x"c0"),
  2568 => (x"c4",x"01",x"a9",x"c0"),
  2569 => (x"c2",x"4a",x"c0",x"87"),
  2570 => (x"72",x"4a",x"c1",x"87"),
  2571 => (x"0e",x"4f",x"26",x"48"),
  2572 => (x"5d",x"5c",x"5b",x"5e"),
  2573 => (x"4d",x"71",x"1e",x"0e"),
  2574 => (x"75",x"4b",x"d4",x"ff"),
  2575 => (x"fa",x"cd",x"c3",x"1e"),
  2576 => (x"c2",x"c0",x"fe",x"49"),
  2577 => (x"70",x"86",x"c4",x"87"),
  2578 => (x"c3",x"02",x"6e",x"7e"),
  2579 => (x"ce",x"c3",x"87",x"ff"),
  2580 => (x"75",x"4c",x"bf",x"c2"),
  2581 => (x"f0",x"d9",x"fe",x"49"),
  2582 => (x"05",x"a8",x"de",x"87"),
  2583 => (x"75",x"87",x"eb",x"c0"),
  2584 => (x"f6",x"d0",x"ff",x"49"),
  2585 => (x"02",x"98",x"70",x"87"),
  2586 => (x"cc",x"c3",x"87",x"db"),
  2587 => (x"c0",x"1e",x"bf",x"fd"),
  2588 => (x"ce",x"ff",x"49",x"e1"),
  2589 => (x"86",x"c4",x"87",x"c9"),
  2590 => (x"48",x"e7",x"e5",x"c2"),
  2591 => (x"cd",x"c3",x"50",x"c0"),
  2592 => (x"ea",x"fe",x"49",x"c9"),
  2593 => (x"c3",x"48",x"c1",x"87"),
  2594 => (x"d0",x"ff",x"87",x"c5"),
  2595 => (x"78",x"c5",x"c8",x"48"),
  2596 => (x"c0",x"7b",x"d6",x"c1"),
  2597 => (x"bf",x"97",x"6e",x"4a"),
  2598 => (x"c1",x"48",x"6e",x"7b"),
  2599 => (x"c1",x"7e",x"70",x"80"),
  2600 => (x"b7",x"e0",x"c0",x"82"),
  2601 => (x"ec",x"ff",x"04",x"aa"),
  2602 => (x"48",x"d0",x"ff",x"87"),
  2603 => (x"c5",x"c8",x"78",x"c4"),
  2604 => (x"7b",x"d3",x"c1",x"78"),
  2605 => (x"78",x"c4",x"7b",x"c1"),
  2606 => (x"c1",x"02",x"9c",x"74"),
  2607 => (x"fb",x"c2",x"87",x"fd"),
  2608 => (x"c0",x"c8",x"7e",x"f6"),
  2609 => (x"b7",x"c0",x"8c",x"4d"),
  2610 => (x"87",x"c6",x"03",x"ac"),
  2611 => (x"4d",x"a4",x"c0",x"c8"),
  2612 => (x"c8",x"c3",x"4c",x"c0"),
  2613 => (x"49",x"bf",x"97",x"e7"),
  2614 => (x"d2",x"02",x"99",x"d0"),
  2615 => (x"c3",x"1e",x"c0",x"87"),
  2616 => (x"fe",x"49",x"fa",x"cd"),
  2617 => (x"c4",x"87",x"fc",x"c0"),
  2618 => (x"4a",x"49",x"70",x"86"),
  2619 => (x"c2",x"87",x"ef",x"c0"),
  2620 => (x"c3",x"1e",x"f6",x"fb"),
  2621 => (x"fe",x"49",x"fa",x"cd"),
  2622 => (x"c4",x"87",x"e8",x"c0"),
  2623 => (x"4a",x"49",x"70",x"86"),
  2624 => (x"c8",x"48",x"d0",x"ff"),
  2625 => (x"d4",x"c1",x"78",x"c5"),
  2626 => (x"bf",x"97",x"6e",x"7b"),
  2627 => (x"c1",x"48",x"6e",x"7b"),
  2628 => (x"c1",x"7e",x"70",x"80"),
  2629 => (x"f0",x"ff",x"05",x"8d"),
  2630 => (x"48",x"d0",x"ff",x"87"),
  2631 => (x"9a",x"72",x"78",x"c4"),
  2632 => (x"87",x"c5",x"c0",x"05"),
  2633 => (x"e6",x"c0",x"48",x"c0"),
  2634 => (x"c3",x"1e",x"c1",x"87"),
  2635 => (x"fd",x"49",x"fa",x"cd"),
  2636 => (x"c4",x"87",x"cf",x"fe"),
  2637 => (x"05",x"9c",x"74",x"86"),
  2638 => (x"ff",x"87",x"c3",x"fe"),
  2639 => (x"c5",x"c8",x"48",x"d0"),
  2640 => (x"7b",x"d3",x"c1",x"78"),
  2641 => (x"78",x"c4",x"7b",x"c0"),
  2642 => (x"c2",x"c0",x"48",x"c1"),
  2643 => (x"26",x"48",x"c0",x"87"),
  2644 => (x"4c",x"26",x"4d",x"26"),
  2645 => (x"4f",x"26",x"4b",x"26"),
  2646 => (x"c4",x"4a",x"71",x"1e"),
  2647 => (x"87",x"c5",x"05",x"66"),
  2648 => (x"ca",x"fb",x"49",x"72"),
  2649 => (x"00",x"4f",x"26",x"87"),
  2650 => (x"f6",x"e6",x"c2",x"1e"),
  2651 => (x"b9",x"c1",x"49",x"bf"),
  2652 => (x"59",x"fa",x"e6",x"c2"),
  2653 => (x"c3",x"48",x"d4",x"ff"),
  2654 => (x"d0",x"ff",x"78",x"ff"),
  2655 => (x"78",x"e1",x"c8",x"48"),
  2656 => (x"c1",x"48",x"d4",x"ff"),
  2657 => (x"71",x"31",x"c4",x"78"),
  2658 => (x"48",x"d0",x"ff",x"78"),
  2659 => (x"26",x"78",x"e0",x"c0"),
  2660 => (x"e6",x"c2",x"1e",x"4f"),
  2661 => (x"cd",x"c3",x"1e",x"ea"),
  2662 => (x"fa",x"fd",x"49",x"fa"),
  2663 => (x"86",x"c4",x"87",x"e9"),
  2664 => (x"c3",x"02",x"98",x"70"),
  2665 => (x"87",x"c0",x"ff",x"87"),
  2666 => (x"35",x"31",x"4f",x"26"),
  2667 => (x"20",x"5a",x"48",x"4b"),
  2668 => (x"46",x"43",x"20",x"20"),
  2669 => (x"00",x"00",x"00",x"47"),
  2670 => (x"fe",x"1e",x"00",x"00"),
  2671 => (x"c4",x"87",x"f8",x"fd"),
  2672 => (x"c0",x"c2",x"49",x"66"),
  2673 => (x"87",x"cd",x"02",x"99"),
  2674 => (x"c3",x"1e",x"e0",x"c3"),
  2675 => (x"fe",x"49",x"d3",x"cc"),
  2676 => (x"c4",x"87",x"c7",x"ff"),
  2677 => (x"49",x"66",x"c4",x"86"),
  2678 => (x"02",x"99",x"c0",x"c4"),
  2679 => (x"f0",x"c3",x"87",x"cd"),
  2680 => (x"d3",x"cc",x"c3",x"1e"),
  2681 => (x"f1",x"fe",x"fe",x"49"),
  2682 => (x"c4",x"86",x"c4",x"87"),
  2683 => (x"ff",x"c1",x"49",x"66"),
  2684 => (x"c3",x"1e",x"71",x"99"),
  2685 => (x"fe",x"49",x"d3",x"cc"),
  2686 => (x"fe",x"87",x"df",x"fe"),
  2687 => (x"26",x"87",x"f0",x"fc"),
  2688 => (x"5e",x"0e",x"4f",x"26"),
  2689 => (x"0e",x"5d",x"5c",x"5b"),
  2690 => (x"c0",x"86",x"d8",x"ff"),
  2691 => (x"d2",x"ce",x"c3",x"7e"),
  2692 => (x"81",x"c2",x"49",x"bf"),
  2693 => (x"1e",x"72",x"1e",x"71"),
  2694 => (x"db",x"fd",x"4a",x"c6"),
  2695 => (x"48",x"71",x"87",x"e8"),
  2696 => (x"49",x"26",x"4a",x"26"),
  2697 => (x"c3",x"58",x"a6",x"c8"),
  2698 => (x"49",x"bf",x"d2",x"ce"),
  2699 => (x"1e",x"71",x"81",x"c4"),
  2700 => (x"4a",x"c6",x"1e",x"72"),
  2701 => (x"87",x"ce",x"db",x"fd"),
  2702 => (x"4a",x"26",x"48",x"71"),
  2703 => (x"a6",x"cc",x"49",x"26"),
  2704 => (x"d3",x"f3",x"c2",x"58"),
  2705 => (x"cd",x"f7",x"49",x"bf"),
  2706 => (x"02",x"98",x"70",x"87"),
  2707 => (x"c0",x"87",x"f9",x"c9"),
  2708 => (x"f5",x"f6",x"49",x"e0"),
  2709 => (x"c2",x"49",x"70",x"87"),
  2710 => (x"c0",x"59",x"d7",x"f3"),
  2711 => (x"c4",x"49",x"74",x"4c"),
  2712 => (x"81",x"d0",x"fe",x"91"),
  2713 => (x"49",x"74",x"4a",x"69"),
  2714 => (x"bf",x"d2",x"ce",x"c3"),
  2715 => (x"c3",x"91",x"c4",x"81"),
  2716 => (x"72",x"81",x"de",x"ce"),
  2717 => (x"d2",x"02",x"9a",x"79"),
  2718 => (x"c1",x"49",x"72",x"87"),
  2719 => (x"6e",x"9a",x"71",x"89"),
  2720 => (x"70",x"80",x"c1",x"48"),
  2721 => (x"05",x"9a",x"72",x"7e"),
  2722 => (x"c1",x"87",x"ee",x"ff"),
  2723 => (x"ac",x"b7",x"c2",x"84"),
  2724 => (x"87",x"c9",x"ff",x"04"),
  2725 => (x"fc",x"c0",x"48",x"6e"),
  2726 => (x"c8",x"04",x"a8",x"b7"),
  2727 => (x"4c",x"c0",x"87",x"ea"),
  2728 => (x"66",x"c4",x"4a",x"74"),
  2729 => (x"c3",x"92",x"c4",x"82"),
  2730 => (x"74",x"82",x"de",x"ce"),
  2731 => (x"81",x"66",x"c8",x"49"),
  2732 => (x"ce",x"c3",x"91",x"c4"),
  2733 => (x"4a",x"6a",x"81",x"de"),
  2734 => (x"b9",x"72",x"49",x"69"),
  2735 => (x"ce",x"c3",x"4b",x"74"),
  2736 => (x"c4",x"83",x"bf",x"d2"),
  2737 => (x"de",x"ce",x"c3",x"93"),
  2738 => (x"72",x"ba",x"6b",x"83"),
  2739 => (x"d4",x"98",x"71",x"48"),
  2740 => (x"49",x"74",x"58",x"a6"),
  2741 => (x"bf",x"d2",x"ce",x"c3"),
  2742 => (x"c3",x"91",x"c4",x"81"),
  2743 => (x"69",x"81",x"de",x"ce"),
  2744 => (x"48",x"a6",x"d4",x"7e"),
  2745 => (x"a6",x"d0",x"78",x"c0"),
  2746 => (x"4c",x"ff",x"c3",x"5c"),
  2747 => (x"df",x"49",x"66",x"d0"),
  2748 => (x"e2",x"c6",x"02",x"29"),
  2749 => (x"4a",x"66",x"cc",x"87"),
  2750 => (x"d4",x"92",x"e0",x"c0"),
  2751 => (x"ff",x"c0",x"82",x"66"),
  2752 => (x"70",x"88",x"72",x"48"),
  2753 => (x"48",x"a6",x"d8",x"4a"),
  2754 => (x"80",x"c4",x"78",x"c0"),
  2755 => (x"49",x"6e",x"78",x"c0"),
  2756 => (x"e4",x"c0",x"29",x"df"),
  2757 => (x"ce",x"c3",x"59",x"a6"),
  2758 => (x"78",x"c1",x"48",x"ce"),
  2759 => (x"31",x"c3",x"49",x"72"),
  2760 => (x"b1",x"72",x"2a",x"b7"),
  2761 => (x"c4",x"99",x"ff",x"c0"),
  2762 => (x"ce",x"f7",x"c2",x"91"),
  2763 => (x"6d",x"85",x"71",x"4d"),
  2764 => (x"c0",x"c4",x"49",x"4b"),
  2765 => (x"d7",x"02",x"99",x"c0"),
  2766 => (x"66",x"e0",x"c0",x"87"),
  2767 => (x"87",x"c7",x"c0",x"02"),
  2768 => (x"78",x"c0",x"80",x"c8"),
  2769 => (x"c3",x"87",x"d0",x"c5"),
  2770 => (x"c1",x"48",x"d6",x"ce"),
  2771 => (x"87",x"c7",x"c5",x"78"),
  2772 => (x"02",x"66",x"e0",x"c0"),
  2773 => (x"49",x"73",x"87",x"d8"),
  2774 => (x"99",x"c0",x"c0",x"c2"),
  2775 => (x"87",x"c3",x"c0",x"02"),
  2776 => (x"6d",x"2b",x"b7",x"d0"),
  2777 => (x"ff",x"ff",x"fd",x"48"),
  2778 => (x"c0",x"7d",x"70",x"98"),
  2779 => (x"ce",x"c3",x"87",x"fa"),
  2780 => (x"c0",x"02",x"bf",x"d6"),
  2781 => (x"48",x"73",x"87",x"f2"),
  2782 => (x"c0",x"28",x"b7",x"d0"),
  2783 => (x"70",x"58",x"a6",x"e8"),
  2784 => (x"e3",x"c0",x"02",x"98"),
  2785 => (x"da",x"ce",x"c3",x"87"),
  2786 => (x"e0",x"c0",x"49",x"bf"),
  2787 => (x"c0",x"02",x"99",x"c0"),
  2788 => (x"49",x"70",x"87",x"ca"),
  2789 => (x"99",x"c0",x"e0",x"c0"),
  2790 => (x"87",x"cc",x"c0",x"02"),
  2791 => (x"c0",x"c2",x"48",x"6d"),
  2792 => (x"7d",x"70",x"b0",x"c0"),
  2793 => (x"4b",x"66",x"e4",x"c0"),
  2794 => (x"c0",x"c8",x"49",x"73"),
  2795 => (x"c2",x"02",x"99",x"c0"),
  2796 => (x"ce",x"c3",x"87",x"c5"),
  2797 => (x"cc",x"4a",x"bf",x"da"),
  2798 => (x"c0",x"02",x"9a",x"c0"),
  2799 => (x"c0",x"c4",x"87",x"cf"),
  2800 => (x"d7",x"c0",x"02",x"8a"),
  2801 => (x"c0",x"02",x"8a",x"87"),
  2802 => (x"dc",x"c1",x"87",x"f8"),
  2803 => (x"74",x"49",x"73",x"87"),
  2804 => (x"c2",x"91",x"c2",x"99"),
  2805 => (x"11",x"81",x"c2",x"f7"),
  2806 => (x"87",x"db",x"c1",x"4b"),
  2807 => (x"99",x"74",x"49",x"73"),
  2808 => (x"f7",x"c2",x"91",x"c2"),
  2809 => (x"81",x"c1",x"81",x"c2"),
  2810 => (x"e0",x"c0",x"4b",x"11"),
  2811 => (x"c8",x"c0",x"02",x"66"),
  2812 => (x"48",x"a6",x"dc",x"87"),
  2813 => (x"fe",x"c0",x"78",x"d2"),
  2814 => (x"48",x"a6",x"d8",x"87"),
  2815 => (x"c0",x"78",x"d2",x"c4"),
  2816 => (x"49",x"73",x"87",x"f5"),
  2817 => (x"91",x"c2",x"99",x"74"),
  2818 => (x"81",x"c2",x"f7",x"c2"),
  2819 => (x"4b",x"11",x"81",x"c1"),
  2820 => (x"02",x"66",x"e0",x"c0"),
  2821 => (x"dc",x"87",x"c9",x"c0"),
  2822 => (x"d9",x"c1",x"48",x"a6"),
  2823 => (x"87",x"d7",x"c0",x"78"),
  2824 => (x"c5",x"48",x"a6",x"d8"),
  2825 => (x"ce",x"c0",x"78",x"d9"),
  2826 => (x"74",x"49",x"73",x"87"),
  2827 => (x"c2",x"91",x"c2",x"99"),
  2828 => (x"c1",x"81",x"c2",x"f7"),
  2829 => (x"c0",x"4b",x"11",x"81"),
  2830 => (x"c0",x"02",x"66",x"e0"),
  2831 => (x"49",x"73",x"87",x"db"),
  2832 => (x"fc",x"c7",x"b9",x"ff"),
  2833 => (x"48",x"71",x"99",x"c0"),
  2834 => (x"bf",x"da",x"ce",x"c3"),
  2835 => (x"de",x"ce",x"c3",x"98"),
  2836 => (x"c4",x"9b",x"74",x"58"),
  2837 => (x"d3",x"c0",x"b3",x"c0"),
  2838 => (x"c7",x"49",x"73",x"87"),
  2839 => (x"71",x"99",x"c0",x"fc"),
  2840 => (x"da",x"ce",x"c3",x"48"),
  2841 => (x"ce",x"c3",x"b0",x"bf"),
  2842 => (x"9b",x"74",x"58",x"de"),
  2843 => (x"c0",x"02",x"66",x"d8"),
  2844 => (x"c3",x"1e",x"87",x"ca"),
  2845 => (x"f5",x"49",x"ce",x"ce"),
  2846 => (x"86",x"c4",x"87",x"c0"),
  2847 => (x"ce",x"c3",x"1e",x"73"),
  2848 => (x"f5",x"f4",x"49",x"ce"),
  2849 => (x"dc",x"86",x"c4",x"87"),
  2850 => (x"ca",x"c0",x"02",x"66"),
  2851 => (x"ce",x"c3",x"1e",x"87"),
  2852 => (x"e5",x"f4",x"49",x"ce"),
  2853 => (x"d0",x"86",x"c4",x"87"),
  2854 => (x"30",x"c1",x"48",x"66"),
  2855 => (x"6e",x"58",x"a6",x"d4"),
  2856 => (x"70",x"30",x"c1",x"48"),
  2857 => (x"48",x"66",x"d4",x"7e"),
  2858 => (x"a6",x"d8",x"80",x"c1"),
  2859 => (x"b7",x"e0",x"c0",x"58"),
  2860 => (x"f7",x"f8",x"04",x"a8"),
  2861 => (x"4c",x"66",x"cc",x"87"),
  2862 => (x"b7",x"c2",x"84",x"c1"),
  2863 => (x"df",x"f7",x"04",x"ac"),
  2864 => (x"d2",x"ce",x"c3",x"87"),
  2865 => (x"78",x"66",x"c4",x"48"),
  2866 => (x"26",x"8e",x"d8",x"ff"),
  2867 => (x"26",x"4c",x"26",x"4d"),
  2868 => (x"00",x"4f",x"26",x"4b"),
  2869 => (x"1e",x"00",x"00",x"00"),
  2870 => (x"49",x"72",x"4a",x"c0"),
  2871 => (x"ce",x"c3",x"91",x"c4"),
  2872 => (x"79",x"ff",x"81",x"de"),
  2873 => (x"b7",x"c6",x"82",x"c1"),
  2874 => (x"87",x"ee",x"04",x"aa"),
  2875 => (x"48",x"d2",x"ce",x"c3"),
  2876 => (x"78",x"40",x"40",x"c0"),
  2877 => (x"73",x"1e",x"4f",x"26"),
  2878 => (x"f4",x"4b",x"71",x"1e"),
  2879 => (x"49",x"73",x"87",x"c4"),
  2880 => (x"87",x"c7",x"f6",x"fe"),
  2881 => (x"0e",x"87",x"c8",x"ff"),
  2882 => (x"0e",x"5c",x"5b",x"5e"),
  2883 => (x"ff",x"4c",x"d4",x"ff"),
  2884 => (x"c5",x"c8",x"4b",x"d0"),
  2885 => (x"7c",x"d5",x"c1",x"7b"),
  2886 => (x"c4",x"7c",x"66",x"cc"),
  2887 => (x"7b",x"c5",x"c8",x"7b"),
  2888 => (x"c1",x"7c",x"d3",x"c1"),
  2889 => (x"c8",x"7b",x"c4",x"7c"),
  2890 => (x"d4",x"c1",x"7b",x"c5"),
  2891 => (x"b7",x"4a",x"c0",x"7c"),
  2892 => (x"87",x"cb",x"06",x"a9"),
  2893 => (x"c1",x"7c",x"ff",x"c3"),
  2894 => (x"aa",x"b7",x"71",x"82"),
  2895 => (x"c4",x"87",x"f5",x"04"),
  2896 => (x"7b",x"c5",x"c8",x"7b"),
  2897 => (x"c0",x"7c",x"d3",x"c1"),
  2898 => (x"fd",x"7b",x"c4",x"7c"),
  2899 => (x"73",x"1e",x"87",x"ff"),
  2900 => (x"49",x"4b",x"71",x"1e"),
  2901 => (x"e2",x"c1",x"91",x"cb"),
  2902 => (x"82",x"71",x"4a",x"ee"),
  2903 => (x"97",x"e5",x"cd",x"c3"),
  2904 => (x"87",x"d3",x"02",x"bf"),
  2905 => (x"11",x"49",x"a2",x"ca"),
  2906 => (x"c1",x"87",x"cc",x"05"),
  2907 => (x"49",x"c0",x"c8",x"1e"),
  2908 => (x"c4",x"87",x"d4",x"fe"),
  2909 => (x"73",x"87",x"cc",x"86"),
  2910 => (x"f7",x"d4",x"fe",x"49"),
  2911 => (x"fe",x"49",x"73",x"87"),
  2912 => (x"fd",x"87",x"f1",x"d4"),
  2913 => (x"73",x"1e",x"87",x"c9"),
  2914 => (x"c2",x"4b",x"c0",x"1e"),
  2915 => (x"ea",x"49",x"e3",x"f6"),
  2916 => (x"98",x"70",x"87",x"dd"),
  2917 => (x"c2",x"87",x"c4",x"05"),
  2918 => (x"fc",x"4b",x"ef",x"f6"),
  2919 => (x"48",x"73",x"87",x"f9"),
  2920 => (x"53",x"87",x"ec",x"fc"),
  2921 => (x"32",x"33",x"49",x"56"),
  2922 => (x"52",x"20",x"20",x"38"),
  2923 => (x"52",x"00",x"4d",x"4f"),
  2924 => (x"6c",x"20",x"4d",x"4f"),
  2925 => (x"69",x"64",x"61",x"6f"),
  2926 => (x"66",x"20",x"67",x"6e"),
  2927 => (x"65",x"6c",x"69",x"61"),
  2928 => (x"eb",x"f4",x"00",x"64"),
  2929 => (x"06",x"05",x"f5",x"f2"),
  2930 => (x"0b",x"03",x"0c",x"04"),
  2931 => (x"00",x"66",x"0a",x"83"),
  2932 => (x"00",x"5a",x"00",x"fc"),
  2933 => (x"80",x"00",x"00",x"da"),
  2934 => (x"80",x"05",x"08",x"94"),
  2935 => (x"80",x"02",x"00",x"78"),
  2936 => (x"80",x"03",x"00",x"01"),
  2937 => (x"80",x"04",x"00",x"09"),
  2938 => (x"80",x"01",x"00",x"00"),
  2939 => (x"00",x"26",x"08",x"91"),
  2940 => (x"00",x"1d",x"00",x"04"),
  2941 => (x"00",x"1c",x"00",x"00"),
  2942 => (x"00",x"25",x"00",x"00"),
  2943 => (x"00",x"1a",x"00",x"0c"),
  2944 => (x"00",x"1b",x"00",x"00"),
  2945 => (x"00",x"24",x"00",x"00"),
  2946 => (x"01",x"12",x"00",x"00"),
  2947 => (x"00",x"2e",x"00",x"00"),
  2948 => (x"00",x"2d",x"00",x"03"),
  2949 => (x"00",x"23",x"00",x"00"),
  2950 => (x"00",x"36",x"00",x"00"),
  2951 => (x"00",x"21",x"00",x"0b"),
  2952 => (x"00",x"2b",x"00",x"00"),
  2953 => (x"00",x"2c",x"00",x"00"),
  2954 => (x"00",x"22",x"00",x"00"),
  2955 => (x"00",x"3d",x"00",x"00"),
  2956 => (x"00",x"35",x"00",x"6c"),
  2957 => (x"00",x"34",x"00",x"00"),
  2958 => (x"00",x"3e",x"00",x"00"),
  2959 => (x"00",x"32",x"00",x"75"),
  2960 => (x"00",x"33",x"00",x"00"),
  2961 => (x"00",x"3c",x"00",x"00"),
  2962 => (x"00",x"2a",x"00",x"6b"),
  2963 => (x"00",x"46",x"00",x"00"),
  2964 => (x"00",x"43",x"00",x"01"),
  2965 => (x"00",x"3b",x"00",x"73"),
  2966 => (x"00",x"45",x"00",x"69"),
  2967 => (x"00",x"3a",x"00",x"09"),
  2968 => (x"00",x"42",x"00",x"70"),
  2969 => (x"00",x"44",x"00",x"72"),
  2970 => (x"00",x"31",x"00",x"74"),
  2971 => (x"00",x"55",x"00",x"00"),
  2972 => (x"00",x"4d",x"00",x"00"),
  2973 => (x"00",x"4b",x"00",x"7c"),
  2974 => (x"00",x"7b",x"00",x"7a"),
  2975 => (x"00",x"49",x"00",x"00"),
  2976 => (x"00",x"4c",x"00",x"71"),
  2977 => (x"00",x"54",x"00",x"84"),
  2978 => (x"00",x"41",x"00",x"77"),
  2979 => (x"00",x"61",x"00",x"00"),
  2980 => (x"00",x"5b",x"00",x"00"),
  2981 => (x"00",x"52",x"00",x"7c"),
  2982 => (x"00",x"f1",x"00",x"00"),
  2983 => (x"02",x"59",x"00",x"00"),
  2984 => (x"00",x"0e",x"00",x"00"),
  2985 => (x"00",x"5d",x"00",x"5d"),
  2986 => (x"00",x"4a",x"00",x"00"),
  2987 => (x"00",x"16",x"00",x"79"),
  2988 => (x"00",x"76",x"00",x"05"),
  2989 => (x"00",x"0d",x"00",x"07"),
  2990 => (x"00",x"1e",x"00",x"0d"),
  2991 => (x"00",x"29",x"00",x"06"),
  2992 => (x"04",x"14",x"00",x"00"),
  2993 => (x"00",x"15",x"00",x"00"),
  2994 => (x"40",x"00",x"00",x"00"),
  2995 => (x"40",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

