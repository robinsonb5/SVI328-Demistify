library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"f8cec387",
    12 => x"86c0c64e",
    13 => x"49f8cec3",
    14 => x"48d0fbc2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087ffe0",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"4a66c41e",
    47 => x"51124871",
    48 => x"2687fb05",
    49 => x"48731e4f",
    50 => x"05a97381",
    51 => x"87f95372",
    52 => x"731e4f26",
    53 => x"029a721e",
    54 => x"c087e7c0",
    55 => x"724bc148",
    56 => x"87d106a9",
    57 => x"c9068272",
    58 => x"72837387",
    59 => x"87f401a9",
    60 => x"b2c187c3",
    61 => x"03a9723a",
    62 => x"07807389",
    63 => x"052b2ac1",
    64 => x"4b2687f3",
    65 => x"751e4f26",
    66 => x"714dc41e",
    67 => x"ff04a1b7",
    68 => x"c381c1b9",
    69 => x"b77207bd",
    70 => x"baff04a2",
    71 => x"bdc182c1",
    72 => x"87eefe07",
    73 => x"ff042dc1",
    74 => x"0780c1b8",
    75 => x"b9ff042d",
    76 => x"260781c1",
    77 => x"1e4f264d",
    78 => x"c348d4ff",
    79 => x"516878ff",
    80 => x"c14866c4",
    81 => x"58a6c888",
    82 => x"eb059870",
    83 => x"1e4f2687",
    84 => x"d4ff1e73",
    85 => x"7bffc34b",
    86 => x"ffc34a6b",
    87 => x"c8496b7b",
    88 => x"c3b17232",
    89 => x"4a6b7bff",
    90 => x"b27131c8",
    91 => x"6b7bffc3",
    92 => x"7232c849",
    93 => x"c44871b1",
    94 => x"264d2687",
    95 => x"264b264c",
    96 => x"5b5e0e4f",
    97 => x"710e5d5c",
    98 => x"4cd4ff4a",
    99 => x"ffc34972",
   100 => x"c27c7199",
   101 => x"05bfd0fb",
   102 => x"66d087c8",
   103 => x"d430c948",
   104 => x"66d058a6",
   105 => x"c329d849",
   106 => x"7c7199ff",
   107 => x"d04966d0",
   108 => x"99ffc329",
   109 => x"66d07c71",
   110 => x"c329c849",
   111 => x"7c7199ff",
   112 => x"c34966d0",
   113 => x"7c7199ff",
   114 => x"29d04972",
   115 => x"7199ffc3",
   116 => x"c94b6c7c",
   117 => x"c34dfff0",
   118 => x"d005abff",
   119 => x"7cffc387",
   120 => x"8dc14b6c",
   121 => x"c387c602",
   122 => x"f002abff",
   123 => x"fe487387",
   124 => x"c01e87c7",
   125 => x"48d4ff49",
   126 => x"c178ffc3",
   127 => x"b7c8c381",
   128 => x"87f104a9",
   129 => x"731e4f26",
   130 => x"c487e71e",
   131 => x"c04bdff8",
   132 => x"f0ffc01e",
   133 => x"fd49f7c1",
   134 => x"86c487e7",
   135 => x"c005a8c1",
   136 => x"d4ff87ea",
   137 => x"78ffc348",
   138 => x"c0c0c0c1",
   139 => x"c01ec0c0",
   140 => x"e9c1f0e1",
   141 => x"87c9fd49",
   142 => x"987086c4",
   143 => x"ff87ca05",
   144 => x"ffc348d4",
   145 => x"cb48c178",
   146 => x"87e6fe87",
   147 => x"fe058bc1",
   148 => x"48c087fd",
   149 => x"1e87e6fc",
   150 => x"d4ff1e73",
   151 => x"78ffc348",
   152 => x"1ec04bd3",
   153 => x"c1f0ffc0",
   154 => x"d4fc49c1",
   155 => x"7086c487",
   156 => x"87ca0598",
   157 => x"c348d4ff",
   158 => x"48c178ff",
   159 => x"f1fd87cb",
   160 => x"058bc187",
   161 => x"c087dbff",
   162 => x"87f1fb48",
   163 => x"5c5b5e0e",
   164 => x"4cd4ff0e",
   165 => x"c687dbfd",
   166 => x"e1c01eea",
   167 => x"49c8c1f0",
   168 => x"c487defb",
   169 => x"02a8c186",
   170 => x"eafe87c8",
   171 => x"c148c087",
   172 => x"dafa87e2",
   173 => x"cf497087",
   174 => x"c699ffff",
   175 => x"c802a9ea",
   176 => x"87d3fe87",
   177 => x"cbc148c0",
   178 => x"7cffc387",
   179 => x"fc4bf1c0",
   180 => x"987087f4",
   181 => x"87ebc002",
   182 => x"ffc01ec0",
   183 => x"49fac1f0",
   184 => x"c487defa",
   185 => x"05987086",
   186 => x"ffc387d9",
   187 => x"c3496c7c",
   188 => x"7c7c7cff",
   189 => x"99c0c17c",
   190 => x"c187c402",
   191 => x"c087d548",
   192 => x"c287d148",
   193 => x"87c405ab",
   194 => x"87c848c0",
   195 => x"fe058bc1",
   196 => x"48c087fd",
   197 => x"1e87e4f9",
   198 => x"fbc21e73",
   199 => x"78c148d0",
   200 => x"d0ff4bc7",
   201 => x"fb78c248",
   202 => x"d0ff87c8",
   203 => x"c078c348",
   204 => x"d0e5c01e",
   205 => x"f949c0c1",
   206 => x"86c487c7",
   207 => x"c105a8c1",
   208 => x"abc24b87",
   209 => x"c087c505",
   210 => x"87f9c048",
   211 => x"ff058bc1",
   212 => x"f7fc87d0",
   213 => x"d4fbc287",
   214 => x"05987058",
   215 => x"1ec187cd",
   216 => x"c1f0ffc0",
   217 => x"d8f849d0",
   218 => x"ff86c487",
   219 => x"ffc348d4",
   220 => x"87fec278",
   221 => x"58d8fbc2",
   222 => x"c248d0ff",
   223 => x"48d4ff78",
   224 => x"c178ffc3",
   225 => x"87f5f748",
   226 => x"4ad4ff1e",
   227 => x"c448d0ff",
   228 => x"ffc378d1",
   229 => x"0589c17a",
   230 => x"4f2687f8",
   231 => x"711e731e",
   232 => x"cdeec54b",
   233 => x"d4ff4adf",
   234 => x"78ffc348",
   235 => x"fec34868",
   236 => x"87c502a8",
   237 => x"ed058ac1",
   238 => x"059a7287",
   239 => x"48c087c5",
   240 => x"7387eac0",
   241 => x"87cc029b",
   242 => x"731e66c8",
   243 => x"87e7f549",
   244 => x"87c686c4",
   245 => x"fe4966c8",
   246 => x"d4ff87ee",
   247 => x"78ffc348",
   248 => x"059b7378",
   249 => x"d0ff87c5",
   250 => x"c178d048",
   251 => x"87cdf648",
   252 => x"711e731e",
   253 => x"ff4bc04a",
   254 => x"ffc348d4",
   255 => x"48d0ff78",
   256 => x"ff78c3c4",
   257 => x"ffc348d4",
   258 => x"c01e7278",
   259 => x"d1c1f0ff",
   260 => x"87edf549",
   261 => x"987086c4",
   262 => x"c887cd05",
   263 => x"66cc1ec0",
   264 => x"87f8fd49",
   265 => x"4b7086c4",
   266 => x"c248d0ff",
   267 => x"f5487378",
   268 => x"5e0e87cb",
   269 => x"0e5d5c5b",
   270 => x"ffc01ec0",
   271 => x"49c9c1f0",
   272 => x"d287fef4",
   273 => x"d8fbc21e",
   274 => x"87d0fd49",
   275 => x"4cc086c8",
   276 => x"b7d284c1",
   277 => x"87f804ac",
   278 => x"97d8fbc2",
   279 => x"c0c349bf",
   280 => x"a9c0c199",
   281 => x"87e7c005",
   282 => x"97dffbc2",
   283 => x"31d049bf",
   284 => x"97e0fbc2",
   285 => x"32c84abf",
   286 => x"fbc2b172",
   287 => x"4abf97e1",
   288 => x"cf4c71b1",
   289 => x"9cffffff",
   290 => x"34ca84c1",
   291 => x"c287e7c1",
   292 => x"bf97e1fb",
   293 => x"c631c149",
   294 => x"e2fbc299",
   295 => x"c74abf97",
   296 => x"b1722ab7",
   297 => x"97ddfbc2",
   298 => x"cf4d4abf",
   299 => x"defbc29d",
   300 => x"c34abf97",
   301 => x"c232ca9a",
   302 => x"bf97dffb",
   303 => x"7333c24b",
   304 => x"e0fbc2b2",
   305 => x"c34bbf97",
   306 => x"b7c69bc0",
   307 => x"c2b2732b",
   308 => x"7148c181",
   309 => x"c1497030",
   310 => x"70307548",
   311 => x"c14c724d",
   312 => x"c8947184",
   313 => x"06adb7c0",
   314 => x"34c187cc",
   315 => x"c0c82db7",
   316 => x"ff01adb7",
   317 => x"487487f4",
   318 => x"0e87fef1",
   319 => x"5d5c5b5e",
   320 => x"c386f80e",
   321 => x"c048fec3",
   322 => x"f6fbc278",
   323 => x"fb49c01e",
   324 => x"86c487de",
   325 => x"c5059870",
   326 => x"c948c087",
   327 => x"4dc087ce",
   328 => x"f6c07ec1",
   329 => x"c249bfef",
   330 => x"714aecfc",
   331 => x"f9ec4bc8",
   332 => x"05987087",
   333 => x"7ec087c2",
   334 => x"bfebf6c0",
   335 => x"c8fdc249",
   336 => x"4bc8714a",
   337 => x"7087e3ec",
   338 => x"87c20598",
   339 => x"026e7ec0",
   340 => x"c387fdc0",
   341 => x"4dbffcc2",
   342 => x"9ff4c3c3",
   343 => x"c5487ebf",
   344 => x"05a8ead6",
   345 => x"c2c387c7",
   346 => x"ce4dbffc",
   347 => x"ca486e87",
   348 => x"02a8d5e9",
   349 => x"48c087c5",
   350 => x"c287f1c7",
   351 => x"751ef6fb",
   352 => x"87ecf949",
   353 => x"987086c4",
   354 => x"c087c505",
   355 => x"87dcc748",
   356 => x"bfebf6c0",
   357 => x"c8fdc249",
   358 => x"4bc8714a",
   359 => x"7087cbeb",
   360 => x"87c80598",
   361 => x"48fec3c3",
   362 => x"87da78c1",
   363 => x"bfeff6c0",
   364 => x"ecfcc249",
   365 => x"4bc8714a",
   366 => x"7087efea",
   367 => x"c5c00298",
   368 => x"c648c087",
   369 => x"c3c387e6",
   370 => x"49bf97f4",
   371 => x"05a9d5c1",
   372 => x"c387cdc0",
   373 => x"bf97f5c3",
   374 => x"a9eac249",
   375 => x"87c5c002",
   376 => x"c7c648c0",
   377 => x"f6fbc287",
   378 => x"487ebf97",
   379 => x"02a8e9c3",
   380 => x"6e87cec0",
   381 => x"a8ebc348",
   382 => x"87c5c002",
   383 => x"ebc548c0",
   384 => x"c1fcc287",
   385 => x"9949bf97",
   386 => x"87ccc005",
   387 => x"97c2fcc2",
   388 => x"a9c249bf",
   389 => x"87c5c002",
   390 => x"cfc548c0",
   391 => x"c3fcc287",
   392 => x"c348bf97",
   393 => x"7058fac3",
   394 => x"88c1484c",
   395 => x"58fec3c3",
   396 => x"97c4fcc2",
   397 => x"817549bf",
   398 => x"97c5fcc2",
   399 => x"32c84abf",
   400 => x"c37ea172",
   401 => x"6e48cbc8",
   402 => x"c6fcc278",
   403 => x"c848bf97",
   404 => x"c3c358a6",
   405 => x"c202bffe",
   406 => x"f6c087d4",
   407 => x"c249bfeb",
   408 => x"714ac8fd",
   409 => x"c1e84bc8",
   410 => x"02987087",
   411 => x"c087c5c0",
   412 => x"87f8c348",
   413 => x"bff6c3c3",
   414 => x"dfc8c34c",
   415 => x"dbfcc25c",
   416 => x"c849bf97",
   417 => x"dafcc231",
   418 => x"a14abf97",
   419 => x"dcfcc249",
   420 => x"d04abf97",
   421 => x"49a17232",
   422 => x"97ddfcc2",
   423 => x"32d84abf",
   424 => x"c449a172",
   425 => x"c8c39166",
   426 => x"c381bfcb",
   427 => x"c259d3c8",
   428 => x"bf97e3fc",
   429 => x"c232c84a",
   430 => x"bf97e2fc",
   431 => x"c24aa24b",
   432 => x"bf97e4fc",
   433 => x"7333d04b",
   434 => x"fcc24aa2",
   435 => x"4bbf97e5",
   436 => x"33d89bcf",
   437 => x"c34aa273",
   438 => x"c35ad7c8",
   439 => x"4abfd3c8",
   440 => x"92748ac2",
   441 => x"48d7c8c3",
   442 => x"c178a172",
   443 => x"fcc287ca",
   444 => x"49bf97c8",
   445 => x"fcc231c8",
   446 => x"4abf97c7",
   447 => x"c4c349a1",
   448 => x"c4c359c6",
   449 => x"c549bfc2",
   450 => x"81ffc731",
   451 => x"c8c329c9",
   452 => x"fcc259df",
   453 => x"4abf97cd",
   454 => x"fcc232c8",
   455 => x"4bbf97cc",
   456 => x"66c44aa2",
   457 => x"c3826e92",
   458 => x"c35adbc8",
   459 => x"c048d3c8",
   460 => x"cfc8c378",
   461 => x"78a17248",
   462 => x"48dfc8c3",
   463 => x"bfd3c8c3",
   464 => x"e3c8c378",
   465 => x"d7c8c348",
   466 => x"c3c378bf",
   467 => x"c002bffe",
   468 => x"487487c9",
   469 => x"7e7030c4",
   470 => x"c387c9c0",
   471 => x"48bfdbc8",
   472 => x"7e7030c4",
   473 => x"48c2c4c3",
   474 => x"48c1786e",
   475 => x"4d268ef8",
   476 => x"4b264c26",
   477 => x"5e0e4f26",
   478 => x"0e5d5c5b",
   479 => x"c3c34a71",
   480 => x"cb02bffe",
   481 => x"c74b7287",
   482 => x"c14c722b",
   483 => x"87c99cff",
   484 => x"2bc84b72",
   485 => x"ffc34c72",
   486 => x"cbc8c39c",
   487 => x"f6c083bf",
   488 => x"02abbfe7",
   489 => x"f6c087d9",
   490 => x"fbc25beb",
   491 => x"49731ef6",
   492 => x"c487fdf0",
   493 => x"05987086",
   494 => x"48c087c5",
   495 => x"c387e6c0",
   496 => x"02bffec3",
   497 => x"497487d2",
   498 => x"fbc291c4",
   499 => x"4d6981f6",
   500 => x"ffffffcf",
   501 => x"87cb9dff",
   502 => x"91c24974",
   503 => x"81f6fbc2",
   504 => x"754d699f",
   505 => x"87c6fe48",
   506 => x"5c5b5e0e",
   507 => x"711e0e5d",
   508 => x"c11ec04d",
   509 => x"87d7cf49",
   510 => x"4c7086c4",
   511 => x"c0c1029c",
   512 => x"c6c4c387",
   513 => x"e149754a",
   514 => x"987087c5",
   515 => x"87f1c002",
   516 => x"49754a74",
   517 => x"ebe14bcb",
   518 => x"02987087",
   519 => x"c087e2c0",
   520 => x"029c741e",
   521 => x"a6c487c7",
   522 => x"c578c048",
   523 => x"48a6c487",
   524 => x"66c478c1",
   525 => x"87d7ce49",
   526 => x"4c7086c4",
   527 => x"c0ff059c",
   528 => x"26487487",
   529 => x"0e87e7fc",
   530 => x"5d5c5b5e",
   531 => x"4b711e0e",
   532 => x"87c5059b",
   533 => x"e5c148c0",
   534 => x"4da3c887",
   535 => x"66d47dc0",
   536 => x"d487c702",
   537 => x"05bf9766",
   538 => x"48c087c5",
   539 => x"d487cfc1",
   540 => x"f3fd4966",
   541 => x"9c4c7087",
   542 => x"87c0c102",
   543 => x"6949a4dc",
   544 => x"49a4da7d",
   545 => x"9f4aa3c4",
   546 => x"c3c37a69",
   547 => x"d202bffe",
   548 => x"49a4d487",
   549 => x"c049699f",
   550 => x"7199ffff",
   551 => x"7030d048",
   552 => x"c087c27e",
   553 => x"48496e7e",
   554 => x"7a70806a",
   555 => x"a3cc7bc0",
   556 => x"d0796a49",
   557 => x"79c049a3",
   558 => x"87c24874",
   559 => x"fa2648c0",
   560 => x"5e0e87ec",
   561 => x"0e5d5c5b",
   562 => x"f6c04c71",
   563 => x"78ff48e7",
   564 => x"c1029c74",
   565 => x"a4c887ca",
   566 => x"c1026949",
   567 => x"66d087c2",
   568 => x"82496c4a",
   569 => x"d05aa6d4",
   570 => x"c3b94d66",
   571 => x"4abffac3",
   572 => x"9972baff",
   573 => x"c0029971",
   574 => x"a4c487e4",
   575 => x"f9496b4b",
   576 => x"7b7087f4",
   577 => x"bff6c3c3",
   578 => x"71816c49",
   579 => x"c3b9757c",
   580 => x"4abffac3",
   581 => x"9972baff",
   582 => x"ff059971",
   583 => x"7c7587dc",
   584 => x"1e87cbf9",
   585 => x"4b711e73",
   586 => x"87c7029b",
   587 => x"6949a3c8",
   588 => x"c087c505",
   589 => x"87ebc048",
   590 => x"bfcfc8c3",
   591 => x"49a3c44a",
   592 => x"89c24969",
   593 => x"bff6c3c3",
   594 => x"4aa27191",
   595 => x"bffac3c3",
   596 => x"71996b49",
   597 => x"66c84aa2",
   598 => x"ea49721e",
   599 => x"86c487d2",
   600 => x"f8484970",
   601 => x"5e0e87cc",
   602 => x"0e5d5c5b",
   603 => x"d44b711e",
   604 => x"2cc94c66",
   605 => x"c1029b73",
   606 => x"a3c887cf",
   607 => x"c1026949",
   608 => x"a3d087c7",
   609 => x"7d66d44d",
   610 => x"bffac3c3",
   611 => x"6bb9ff49",
   612 => x"717e994a",
   613 => x"87cd03ac",
   614 => x"cc7d7bc0",
   615 => x"a3c44aa3",
   616 => x"c2796a49",
   617 => x"748c7287",
   618 => x"87dd029c",
   619 => x"49731e49",
   620 => x"c487cffc",
   621 => x"4966d486",
   622 => x"0299ffc7",
   623 => x"fbc287cb",
   624 => x"49731ef6",
   625 => x"c487dcfd",
   626 => x"e1f62686",
   627 => x"5b5e0e87",
   628 => x"f00e5d5c",
   629 => x"59a6d086",
   630 => x"4b66e4c0",
   631 => x"ca0266cc",
   632 => x"80c84887",
   633 => x"bf6e7e70",
   634 => x"c087c505",
   635 => x"87ecc348",
   636 => x"d04c66cc",
   637 => x"c4497384",
   638 => x"786c48a6",
   639 => x"c48166c4",
   640 => x"78bf6e80",
   641 => x"06a966c8",
   642 => x"c44987c6",
   643 => x"4b718966",
   644 => x"01abb7c0",
   645 => x"c34887c4",
   646 => x"66c487c2",
   647 => x"98ffc748",
   648 => x"026e7e70",
   649 => x"c887c9c1",
   650 => x"896e49c0",
   651 => x"fbc24a71",
   652 => x"856e4df6",
   653 => x"06aab773",
   654 => x"724a87c1",
   655 => x"66c44849",
   656 => x"727c7080",
   657 => x"8ac1498b",
   658 => x"d9029971",
   659 => x"66e0c087",
   660 => x"c0501548",
   661 => x"c14866e0",
   662 => x"a6e4c080",
   663 => x"c1497258",
   664 => x"0599718a",
   665 => x"1ec187e7",
   666 => x"f94966d0",
   667 => x"86c487d4",
   668 => x"06abb7c0",
   669 => x"c087e3c1",
   670 => x"c74d66e0",
   671 => x"06abb7ff",
   672 => x"7587e2c0",
   673 => x"4966d01e",
   674 => x"c887d8fa",
   675 => x"486c85c0",
   676 => x"7080c0c8",
   677 => x"8bc0c87c",
   678 => x"66d41ec1",
   679 => x"87e2f849",
   680 => x"eec086c8",
   681 => x"f6fbc287",
   682 => x"4966d01e",
   683 => x"c487f4f9",
   684 => x"f6fbc286",
   685 => x"4849734a",
   686 => x"7c70806c",
   687 => x"8bc14973",
   688 => x"ce029971",
   689 => x"7d971287",
   690 => x"497385c1",
   691 => x"99718bc1",
   692 => x"c087f205",
   693 => x"fe01abb7",
   694 => x"48c187e1",
   695 => x"cdf28ef0",
   696 => x"5b5e0e87",
   697 => x"710e5d5c",
   698 => x"c7029b4b",
   699 => x"4da3c887",
   700 => x"87c5056d",
   701 => x"fdc048ff",
   702 => x"4ca3d087",
   703 => x"ffc7496c",
   704 => x"87d80599",
   705 => x"87c9026c",
   706 => x"49731ec1",
   707 => x"c487f3f6",
   708 => x"f6fbc286",
   709 => x"f849731e",
   710 => x"86c487c9",
   711 => x"aa6d4a6c",
   712 => x"ff87c404",
   713 => x"c187cf48",
   714 => x"49727ca2",
   715 => x"c299ffc7",
   716 => x"9781f6fb",
   717 => x"f5f04869",
   718 => x"1e731e87",
   719 => x"029b4b71",
   720 => x"c387e4c0",
   721 => x"735be3c8",
   722 => x"c38ac24a",
   723 => x"49bff6c3",
   724 => x"cfc8c392",
   725 => x"807248bf",
   726 => x"58e7c8c3",
   727 => x"30c44871",
   728 => x"58c6c4c3",
   729 => x"c387edc0",
   730 => x"c348dfc8",
   731 => x"78bfd3c8",
   732 => x"48e3c8c3",
   733 => x"bfd7c8c3",
   734 => x"fec3c378",
   735 => x"87c902bf",
   736 => x"bff6c3c3",
   737 => x"c731c449",
   738 => x"dbc8c387",
   739 => x"31c449bf",
   740 => x"59c6c4c3",
   741 => x"0e87dbef",
   742 => x"0e5c5b5e",
   743 => x"4bc04a71",
   744 => x"c0029a72",
   745 => x"a2da87e1",
   746 => x"4b699f49",
   747 => x"bffec3c3",
   748 => x"d487cf02",
   749 => x"699f49a2",
   750 => x"ffc04c49",
   751 => x"34d09cff",
   752 => x"4cc087c2",
   753 => x"73b34974",
   754 => x"87edfd49",
   755 => x"0e87e1ee",
   756 => x"5d5c5b5e",
   757 => x"7186f40e",
   758 => x"727ec04a",
   759 => x"87d8029a",
   760 => x"48f2fbc2",
   761 => x"fbc278c0",
   762 => x"c8c348ea",
   763 => x"c278bfe3",
   764 => x"c348eefb",
   765 => x"78bfdfc8",
   766 => x"48d3c4c3",
   767 => x"c4c350c0",
   768 => x"c249bfc2",
   769 => x"4abff2fb",
   770 => x"c403aa71",
   771 => x"497287c0",
   772 => x"c00599cf",
   773 => x"fbc287e1",
   774 => x"fbc21ef6",
   775 => x"c249bfea",
   776 => x"c148eafb",
   777 => x"ff7178a1",
   778 => x"c487c5df",
   779 => x"e3f6c086",
   780 => x"f6fbc248",
   781 => x"c087cc78",
   782 => x"48bfe3f6",
   783 => x"c080e0c0",
   784 => x"c258e7f6",
   785 => x"48bff2fb",
   786 => x"fbc280c1",
   787 => x"a32758f6",
   788 => x"bf00000d",
   789 => x"9d4dbf97",
   790 => x"87e2c202",
   791 => x"02ade5c3",
   792 => x"c087dbc2",
   793 => x"4bbfe3f6",
   794 => x"1149a3cb",
   795 => x"05accf4c",
   796 => x"7587d2c1",
   797 => x"c199df49",
   798 => x"c391cd89",
   799 => x"c181c6c4",
   800 => x"51124aa3",
   801 => x"124aa3c3",
   802 => x"4aa3c551",
   803 => x"a3c75112",
   804 => x"c951124a",
   805 => x"51124aa3",
   806 => x"124aa3ce",
   807 => x"4aa3d051",
   808 => x"a3d25112",
   809 => x"d451124a",
   810 => x"51124aa3",
   811 => x"124aa3d6",
   812 => x"4aa3d851",
   813 => x"a3dc5112",
   814 => x"de51124a",
   815 => x"51124aa3",
   816 => x"f9c07ec1",
   817 => x"c8497487",
   818 => x"eac00599",
   819 => x"d0497487",
   820 => x"87d00599",
   821 => x"c00266dc",
   822 => x"497387ca",
   823 => x"700f66dc",
   824 => x"87d30298",
   825 => x"c6c0056e",
   826 => x"c6c4c387",
   827 => x"c050c048",
   828 => x"48bfe3f6",
   829 => x"c387e7c2",
   830 => x"c048d3c4",
   831 => x"c4c37e50",
   832 => x"c249bfc2",
   833 => x"4abff2fb",
   834 => x"fc04aa71",
   835 => x"c8c387c0",
   836 => x"c005bfe3",
   837 => x"c3c387c8",
   838 => x"c102bffe",
   839 => x"f6c087fe",
   840 => x"78ff48e7",
   841 => x"bfeefbc2",
   842 => x"87cae949",
   843 => x"fbc24970",
   844 => x"a6c459f2",
   845 => x"eefbc248",
   846 => x"c3c378bf",
   847 => x"c002bffe",
   848 => x"66c487d8",
   849 => x"ffffcf49",
   850 => x"a999f8ff",
   851 => x"87c5c002",
   852 => x"e1c04dc0",
   853 => x"c04dc187",
   854 => x"66c487dc",
   855 => x"f8ffcf49",
   856 => x"c002a999",
   857 => x"a6c887c8",
   858 => x"c078c048",
   859 => x"a6c887c5",
   860 => x"c878c148",
   861 => x"9d754d66",
   862 => x"87e0c005",
   863 => x"c24966c4",
   864 => x"f6c3c389",
   865 => x"c3914abf",
   866 => x"4abfcfc8",
   867 => x"48eafbc2",
   868 => x"c278a172",
   869 => x"c048f2fb",
   870 => x"87e2f978",
   871 => x"8ef448c0",
   872 => x"0087cbe7",
   873 => x"ff000000",
   874 => x"b3ffffff",
   875 => x"bc00000d",
   876 => x"4600000d",
   877 => x"32335441",
   878 => x"00202020",
   879 => x"31544146",
   880 => x"20202036",
   881 => x"c8c31e00",
   882 => x"dd48bfe8",
   883 => x"87c905a8",
   884 => x"87e8fdc0",
   885 => x"c84a4970",
   886 => x"48d4ff87",
   887 => x"6878ffc3",
   888 => x"2648724a",
   889 => x"c8c31e4f",
   890 => x"dd48bfe8",
   891 => x"87c605a8",
   892 => x"87f4fcc0",
   893 => x"d4ff87d9",
   894 => x"78ffc348",
   895 => x"c848d0ff",
   896 => x"d4ff78e1",
   897 => x"c378d448",
   898 => x"ff48e7c8",
   899 => x"2650bfd4",
   900 => x"d0ff1e4f",
   901 => x"78e0c048",
   902 => x"fe1e4f26",
   903 => x"497087e7",
   904 => x"87c60299",
   905 => x"05a9fbc0",
   906 => x"487187f1",
   907 => x"5e0e4f26",
   908 => x"710e5c5b",
   909 => x"fe4cc04b",
   910 => x"497087cb",
   911 => x"f9c00299",
   912 => x"a9ecc087",
   913 => x"87f2c002",
   914 => x"02a9fbc0",
   915 => x"cc87ebc0",
   916 => x"03acb766",
   917 => x"66d087c7",
   918 => x"7187c202",
   919 => x"02997153",
   920 => x"84c187c2",
   921 => x"7087defd",
   922 => x"cd029949",
   923 => x"a9ecc087",
   924 => x"c087c702",
   925 => x"ff05a9fb",
   926 => x"66d087d5",
   927 => x"c087c302",
   928 => x"ecc07b97",
   929 => x"87c405a9",
   930 => x"87c54a74",
   931 => x"0ac04a74",
   932 => x"c248728a",
   933 => x"264d2687",
   934 => x"264b264c",
   935 => x"e4fc1e4f",
   936 => x"c0497087",
   937 => x"04a9b7f0",
   938 => x"f9c087ca",
   939 => x"c301a9b7",
   940 => x"89f0c087",
   941 => x"a9b7c1c1",
   942 => x"c187ca04",
   943 => x"01a9b7da",
   944 => x"f7c087c3",
   945 => x"26487189",
   946 => x"5b5e0e4f",
   947 => x"4a710e5c",
   948 => x"724cd4ff",
   949 => x"87eac049",
   950 => x"029b4b70",
   951 => x"8bc187c2",
   952 => x"c848d0ff",
   953 => x"d5c178c5",
   954 => x"c649737c",
   955 => x"e7e5c231",
   956 => x"484abf97",
   957 => x"7c70b071",
   958 => x"c448d0ff",
   959 => x"fe487378",
   960 => x"5e0e87d5",
   961 => x"0e5d5c5b",
   962 => x"4c7186f4",
   963 => x"c048a6c4",
   964 => x"7ea4c878",
   965 => x"49bf976e",
   966 => x"05a9c1c1",
   967 => x"a4c987dd",
   968 => x"49699749",
   969 => x"05a9d2c1",
   970 => x"a4ca87d1",
   971 => x"49699749",
   972 => x"05a9c3c1",
   973 => x"48df87c5",
   974 => x"fa87e1c2",
   975 => x"4bc087e7",
   976 => x"97e1ffc0",
   977 => x"a9c049bf",
   978 => x"fb87cf04",
   979 => x"83c187cc",
   980 => x"97e1ffc0",
   981 => x"06ab49bf",
   982 => x"ffc087f1",
   983 => x"02bf97e1",
   984 => x"e0f987cf",
   985 => x"99497087",
   986 => x"c087c602",
   987 => x"f105a9ec",
   988 => x"f94bc087",
   989 => x"4d7087cf",
   990 => x"cc87caf9",
   991 => x"c4f958a6",
   992 => x"c14a7087",
   993 => x"bf976e83",
   994 => x"c702ad49",
   995 => x"adffc087",
   996 => x"87eac005",
   997 => x"9749a4c9",
   998 => x"66c84969",
   999 => x"87c702a9",
  1000 => x"a8ffc048",
  1001 => x"ca87d705",
  1002 => x"699749a4",
  1003 => x"c602aa49",
  1004 => x"aaffc087",
  1005 => x"c487c705",
  1006 => x"78c148a6",
  1007 => x"ecc087d3",
  1008 => x"87c602ad",
  1009 => x"05adfbc0",
  1010 => x"4bc087c7",
  1011 => x"c148a6c4",
  1012 => x"0266c478",
  1013 => x"f887dcfe",
  1014 => x"487387f7",
  1015 => x"f4fa8ef4",
  1016 => x"5e0e0087",
  1017 => x"0e5d5c5b",
  1018 => x"c04b711e",
  1019 => x"04ab4d4c",
  1020 => x"c087e8c0",
  1021 => x"751ec2fc",
  1022 => x"87c4029d",
  1023 => x"87c24ac0",
  1024 => x"49724ac1",
  1025 => x"c487c8ef",
  1026 => x"c17e7086",
  1027 => x"c2056e84",
  1028 => x"c14c7387",
  1029 => x"06ac7385",
  1030 => x"6e87d8ff",
  1031 => x"4d262648",
  1032 => x"4b264c26",
  1033 => x"5e0e4f26",
  1034 => x"0e5d5c5b",
  1035 => x"494c711e",
  1036 => x"c9c391de",
  1037 => x"85714dc1",
  1038 => x"c1026d97",
  1039 => x"c8c387dd",
  1040 => x"744abfec",
  1041 => x"fe497282",
  1042 => x"7e7087d8",
  1043 => x"f3c0026e",
  1044 => x"f4c8c387",
  1045 => x"cb4a6e4b",
  1046 => x"cbc1ff49",
  1047 => x"cb4b7487",
  1048 => x"eee2c193",
  1049 => x"c183c483",
  1050 => x"747bdfc2",
  1051 => x"d6ccc149",
  1052 => x"c37b7587",
  1053 => x"bf97c0c9",
  1054 => x"c8c31e49",
  1055 => x"e3c149f4",
  1056 => x"86c487d6",
  1057 => x"cbc14974",
  1058 => x"49c087fd",
  1059 => x"87dccdc1",
  1060 => x"48e8c8c3",
  1061 => x"49c178c0",
  1062 => x"2687fedc",
  1063 => x"4c87fffd",
  1064 => x"6964616f",
  1065 => x"2e2e676e",
  1066 => x"5e0e002e",
  1067 => x"710e5c5b",
  1068 => x"c8c34a4b",
  1069 => x"7282bfec",
  1070 => x"87e6fc49",
  1071 => x"029c4c70",
  1072 => x"eb4987c4",
  1073 => x"c8c387d1",
  1074 => x"78c048ec",
  1075 => x"c8dc49c1",
  1076 => x"87ccfd87",
  1077 => x"5c5b5e0e",
  1078 => x"86f40e5d",
  1079 => x"4df6fbc2",
  1080 => x"a6c44cc0",
  1081 => x"c378c048",
  1082 => x"49bfecc8",
  1083 => x"c106a9c0",
  1084 => x"fbc287c1",
  1085 => x"029848f6",
  1086 => x"c087f8c0",
  1087 => x"c81ec2fc",
  1088 => x"87c70266",
  1089 => x"c048a6c4",
  1090 => x"c487c578",
  1091 => x"78c148a6",
  1092 => x"ea4966c4",
  1093 => x"86c487f9",
  1094 => x"84c14d70",
  1095 => x"c14866c4",
  1096 => x"58a6c880",
  1097 => x"bfecc8c3",
  1098 => x"c603ac49",
  1099 => x"059d7587",
  1100 => x"c087c8ff",
  1101 => x"029d754c",
  1102 => x"c087e0c3",
  1103 => x"c81ec2fc",
  1104 => x"87c70266",
  1105 => x"c048a6cc",
  1106 => x"cc87c578",
  1107 => x"78c148a6",
  1108 => x"e94966cc",
  1109 => x"86c487f9",
  1110 => x"026e7e70",
  1111 => x"6e87e9c2",
  1112 => x"9781cb49",
  1113 => x"99d04969",
  1114 => x"87d6c102",
  1115 => x"4aeac2c1",
  1116 => x"91cb4974",
  1117 => x"81eee2c1",
  1118 => x"81c87972",
  1119 => x"7451ffc3",
  1120 => x"c391de49",
  1121 => x"714dc1c9",
  1122 => x"97c1c285",
  1123 => x"49a5c17d",
  1124 => x"c351e0c0",
  1125 => x"bf97c6c4",
  1126 => x"c187d202",
  1127 => x"4ba5c284",
  1128 => x"4ac6c4c3",
  1129 => x"fbfe49db",
  1130 => x"dbc187fe",
  1131 => x"49a5cd87",
  1132 => x"84c151c0",
  1133 => x"6e4ba5c2",
  1134 => x"fe49cb4a",
  1135 => x"c187e9fb",
  1136 => x"c0c187c6",
  1137 => x"49744ae6",
  1138 => x"e2c191cb",
  1139 => x"797281ee",
  1140 => x"97c6c4c3",
  1141 => x"87d802bf",
  1142 => x"91de4974",
  1143 => x"c9c384c1",
  1144 => x"83714bc1",
  1145 => x"4ac6c4c3",
  1146 => x"fafe49dd",
  1147 => x"87d887fa",
  1148 => x"93de4b74",
  1149 => x"83c1c9c3",
  1150 => x"c049a3cb",
  1151 => x"7384c151",
  1152 => x"49cb4a6e",
  1153 => x"87e0fafe",
  1154 => x"c14866c4",
  1155 => x"58a6c880",
  1156 => x"c003acc7",
  1157 => x"056e87c5",
  1158 => x"7487e0fc",
  1159 => x"f78ef448",
  1160 => x"731e87fc",
  1161 => x"494b711e",
  1162 => x"e2c191cb",
  1163 => x"a1c881ee",
  1164 => x"e7e5c24a",
  1165 => x"c9501248",
  1166 => x"ffc04aa1",
  1167 => x"501248e1",
  1168 => x"c9c381ca",
  1169 => x"501148c0",
  1170 => x"97c0c9c3",
  1171 => x"c01e49bf",
  1172 => x"c3dcc149",
  1173 => x"e8c8c387",
  1174 => x"c178de48",
  1175 => x"87f9d549",
  1176 => x"87fef626",
  1177 => x"494a711e",
  1178 => x"e2c191cb",
  1179 => x"81c881ee",
  1180 => x"c8c34811",
  1181 => x"c8c358ec",
  1182 => x"78c048ec",
  1183 => x"d8d549c1",
  1184 => x"1e4f2687",
  1185 => x"c5c149c0",
  1186 => x"4f2687e2",
  1187 => x"0299711e",
  1188 => x"e4c187d2",
  1189 => x"50c048c3",
  1190 => x"c9c180f7",
  1191 => x"e2c140e4",
  1192 => x"87ce78e7",
  1193 => x"48ffe3c1",
  1194 => x"78e0e2c1",
  1195 => x"cac180fc",
  1196 => x"4f2678c3",
  1197 => x"5c5b5e0e",
  1198 => x"4a4c710e",
  1199 => x"e2c192cb",
  1200 => x"a2c882ee",
  1201 => x"4ba2c949",
  1202 => x"1e4b6b97",
  1203 => x"1e496997",
  1204 => x"491282ca",
  1205 => x"87c3e6c0",
  1206 => x"fcd349c0",
  1207 => x"c1497487",
  1208 => x"f887e4c2",
  1209 => x"87f8f48e",
  1210 => x"711e731e",
  1211 => x"4aa3c64b",
  1212 => x"c187db02",
  1213 => x"87d6028a",
  1214 => x"dac1028a",
  1215 => x"c0028a87",
  1216 => x"028a87fc",
  1217 => x"8a87e1c0",
  1218 => x"c187cb02",
  1219 => x"49c787db",
  1220 => x"c187d1fd",
  1221 => x"c8c387de",
  1222 => x"c102bfec",
  1223 => x"c14887cb",
  1224 => x"f0c8c388",
  1225 => x"87c1c158",
  1226 => x"bff0c8c3",
  1227 => x"87f9c002",
  1228 => x"bfecc8c3",
  1229 => x"c380c148",
  1230 => x"c058f0c8",
  1231 => x"c8c387eb",
  1232 => x"c649bfec",
  1233 => x"f0c8c389",
  1234 => x"a9b7c059",
  1235 => x"c387da03",
  1236 => x"c048ecc8",
  1237 => x"c387d278",
  1238 => x"02bff0c8",
  1239 => x"c8c387cb",
  1240 => x"c648bfec",
  1241 => x"f0c8c380",
  1242 => x"d149c058",
  1243 => x"497387eb",
  1244 => x"87d3c0c1",
  1245 => x"1e87ebf2",
  1246 => x"4b711e73",
  1247 => x"48e8c8c3",
  1248 => x"49c078dd",
  1249 => x"7387d2d1",
  1250 => x"faffc049",
  1251 => x"87d2f287",
  1252 => x"5c5b5e0e",
  1253 => x"cc4c710e",
  1254 => x"4b741e66",
  1255 => x"e2c193cb",
  1256 => x"a3c483ee",
  1257 => x"fe496a4a",
  1258 => x"c187cdf4",
  1259 => x"c87be2c8",
  1260 => x"66d449a3",
  1261 => x"49a3c951",
  1262 => x"ca5166d8",
  1263 => x"66dc49a3",
  1264 => x"dbf12651",
  1265 => x"5b5e0e87",
  1266 => x"ff0e5d5c",
  1267 => x"a6dc86cc",
  1268 => x"48a6c859",
  1269 => x"80c478c0",
  1270 => x"7866c8c1",
  1271 => x"78c180c4",
  1272 => x"78c180c4",
  1273 => x"48f0c8c3",
  1274 => x"c8c378c1",
  1275 => x"de48bfe8",
  1276 => x"87cb05a8",
  1277 => x"7087ddf3",
  1278 => x"59a6cc49",
  1279 => x"e787d6ce",
  1280 => x"d5e887e3",
  1281 => x"87fde687",
  1282 => x"fbc04c70",
  1283 => x"d8c102ac",
  1284 => x"0566d887",
  1285 => x"c087cac1",
  1286 => x"1ec11e1e",
  1287 => x"1ed1e4c1",
  1288 => x"ebfd49c0",
  1289 => x"c086d087",
  1290 => x"d902acfb",
  1291 => x"66c4c187",
  1292 => x"6a82c44a",
  1293 => x"7481c749",
  1294 => x"d81ec151",
  1295 => x"c8496a1e",
  1296 => x"87eae781",
  1297 => x"c8c186c8",
  1298 => x"a8c04866",
  1299 => x"c887c701",
  1300 => x"78c148a6",
  1301 => x"c8c187ce",
  1302 => x"88c14866",
  1303 => x"c358a6d0",
  1304 => x"87f6e687",
  1305 => x"c248a6d0",
  1306 => x"029c7478",
  1307 => x"c887e2cc",
  1308 => x"ccc14866",
  1309 => x"cc03a866",
  1310 => x"a6dc87d7",
  1311 => x"e578c048",
  1312 => x"4c7087c3",
  1313 => x"dd4866d8",
  1314 => x"87c605a8",
  1315 => x"d848a6dc",
  1316 => x"d0c17866",
  1317 => x"e8c005ac",
  1318 => x"87e9e487",
  1319 => x"7087e6e4",
  1320 => x"acecc04c",
  1321 => x"e587c505",
  1322 => x"4c7087f0",
  1323 => x"05acd0c1",
  1324 => x"66d487c8",
  1325 => x"d880c148",
  1326 => x"d0c158a6",
  1327 => x"d8ff02ac",
  1328 => x"a6e0c087",
  1329 => x"7866d848",
  1330 => x"c04866dc",
  1331 => x"05a866e0",
  1332 => x"c487d0ca",
  1333 => x"f0c048a6",
  1334 => x"80e0c078",
  1335 => x"c47866d0",
  1336 => x"c478c080",
  1337 => x"7478c080",
  1338 => x"8dfbc04d",
  1339 => x"87ccc902",
  1340 => x"db028dc9",
  1341 => x"028dc287",
  1342 => x"c987cdc1",
  1343 => x"d1c4028d",
  1344 => x"028dc487",
  1345 => x"c187c6c1",
  1346 => x"c5c4028d",
  1347 => x"87e6c887",
  1348 => x"cb4966c8",
  1349 => x"66c4c191",
  1350 => x"4aa1c481",
  1351 => x"1e717e6a",
  1352 => x"48ccdfc1",
  1353 => x"cc4966c4",
  1354 => x"41204aa1",
  1355 => x"ff05aa71",
  1356 => x"511087f8",
  1357 => x"cdc14926",
  1358 => x"dde379f7",
  1359 => x"c04c7087",
  1360 => x"c148a6ec",
  1361 => x"87f4c778",
  1362 => x"c048a6c4",
  1363 => x"4866d078",
  1364 => x"a6d480c1",
  1365 => x"87ede158",
  1366 => x"ecc04c70",
  1367 => x"87d402ac",
  1368 => x"c00266c4",
  1369 => x"a6c887c5",
  1370 => x"7487c95c",
  1371 => x"88f0c048",
  1372 => x"58a6e8c0",
  1373 => x"02acecc0",
  1374 => x"c8e187cc",
  1375 => x"c04c7087",
  1376 => x"ff05acec",
  1377 => x"66c487f4",
  1378 => x"4966d81e",
  1379 => x"66ecc01e",
  1380 => x"d1e4c11e",
  1381 => x"4966d81e",
  1382 => x"c087f5f7",
  1383 => x"c01eca1e",
  1384 => x"cb4966e0",
  1385 => x"66dcc191",
  1386 => x"48a6d881",
  1387 => x"d878a1c4",
  1388 => x"e149bf66",
  1389 => x"86d887f8",
  1390 => x"06a8b7c0",
  1391 => x"c187cac1",
  1392 => x"c81ede1e",
  1393 => x"e149bf66",
  1394 => x"86c887e4",
  1395 => x"c0484970",
  1396 => x"e8c08808",
  1397 => x"b7c058a6",
  1398 => x"ecc006a8",
  1399 => x"66e4c087",
  1400 => x"a8b7dd48",
  1401 => x"87e1c003",
  1402 => x"c049bf6e",
  1403 => x"c08166e4",
  1404 => x"e4c051e0",
  1405 => x"81c14966",
  1406 => x"c281bf6e",
  1407 => x"e4c051c1",
  1408 => x"81c24966",
  1409 => x"c081bf6e",
  1410 => x"a6ecc051",
  1411 => x"c478c148",
  1412 => x"c8e287ea",
  1413 => x"a6e8c087",
  1414 => x"87c1e258",
  1415 => x"58a6f0c0",
  1416 => x"05a8ecc0",
  1417 => x"a687c9c0",
  1418 => x"66e4c048",
  1419 => x"87c4c078",
  1420 => x"87d1deff",
  1421 => x"cb4966c8",
  1422 => x"66c4c191",
  1423 => x"c8807148",
  1424 => x"66c458a6",
  1425 => x"c482c84a",
  1426 => x"81ca4966",
  1427 => x"5166e4c0",
  1428 => x"4966ecc0",
  1429 => x"e4c081c1",
  1430 => x"48c18966",
  1431 => x"49703071",
  1432 => x"977189c1",
  1433 => x"ddccc37a",
  1434 => x"e4c049bf",
  1435 => x"6a972966",
  1436 => x"9871484a",
  1437 => x"58a6f4c0",
  1438 => x"c44966c4",
  1439 => x"c07e6981",
  1440 => x"dc4866e0",
  1441 => x"c002a866",
  1442 => x"a6dc87c8",
  1443 => x"c078c048",
  1444 => x"a6dc87c5",
  1445 => x"dc78c148",
  1446 => x"e0c01e66",
  1447 => x"4966c81e",
  1448 => x"87cadeff",
  1449 => x"4c7086c8",
  1450 => x"06acb7c0",
  1451 => x"6e87d6c1",
  1452 => x"70807448",
  1453 => x"49e0c07e",
  1454 => x"4b6e8974",
  1455 => x"4ac9dfc1",
  1456 => x"e3e7fe71",
  1457 => x"c2486e87",
  1458 => x"c07e7080",
  1459 => x"c14866e8",
  1460 => x"a6ecc080",
  1461 => x"66f0c058",
  1462 => x"7081c149",
  1463 => x"c5c002a9",
  1464 => x"c04dc087",
  1465 => x"4dc187c2",
  1466 => x"a4c21e75",
  1467 => x"48e0c049",
  1468 => x"49708871",
  1469 => x"4966c81e",
  1470 => x"87f2dcff",
  1471 => x"b7c086c8",
  1472 => x"c6ff01a8",
  1473 => x"66e8c087",
  1474 => x"87d3c002",
  1475 => x"c94966c4",
  1476 => x"66e8c081",
  1477 => x"4866c451",
  1478 => x"78f4cac1",
  1479 => x"c487cec0",
  1480 => x"81c94966",
  1481 => x"66c451c2",
  1482 => x"cef5c248",
  1483 => x"a6ecc078",
  1484 => x"c078c148",
  1485 => x"dbff87c6",
  1486 => x"4c7087e0",
  1487 => x"0266ecc0",
  1488 => x"c887f5c0",
  1489 => x"66cc4866",
  1490 => x"cbc004a8",
  1491 => x"4866c887",
  1492 => x"a6cc80c1",
  1493 => x"87e0c058",
  1494 => x"c14866cc",
  1495 => x"58a6d088",
  1496 => x"c187d5c0",
  1497 => x"c005acc6",
  1498 => x"66d087c8",
  1499 => x"d480c148",
  1500 => x"daff58a6",
  1501 => x"4c7087e4",
  1502 => x"c14866d4",
  1503 => x"58a6d880",
  1504 => x"c0029c74",
  1505 => x"66c887cb",
  1506 => x"66ccc148",
  1507 => x"e9f304a8",
  1508 => x"fcd9ff87",
  1509 => x"4866c887",
  1510 => x"c003a8c7",
  1511 => x"c8c387e5",
  1512 => x"78c048f0",
  1513 => x"cb4966c8",
  1514 => x"66c4c191",
  1515 => x"4aa1c481",
  1516 => x"52c04a6a",
  1517 => x"4866c879",
  1518 => x"a6cc80c1",
  1519 => x"04a8c758",
  1520 => x"ff87dbff",
  1521 => x"d5e18ecc",
  1522 => x"00203a87",
  1523 => x"20504944",
  1524 => x"74697753",
  1525 => x"73656863",
  1526 => x"1e731e00",
  1527 => x"029b4b71",
  1528 => x"c8c387c6",
  1529 => x"78c048ec",
  1530 => x"c8c31ec7",
  1531 => x"1e49bfec",
  1532 => x"1eeee2c1",
  1533 => x"bfe8c8c3",
  1534 => x"87c9ef49",
  1535 => x"c8c386cc",
  1536 => x"ea49bfe8",
  1537 => x"9b7387c6",
  1538 => x"c187c802",
  1539 => x"c049eee2",
  1540 => x"e087c6ef",
  1541 => x"c71e87cc",
  1542 => x"49c187d6",
  1543 => x"fe87fafe",
  1544 => x"7087f4eb",
  1545 => x"87cd0298",
  1546 => x"87cff3fe",
  1547 => x"c4029870",
  1548 => x"c24ac187",
  1549 => x"724ac087",
  1550 => x"87ce059a",
  1551 => x"e1c11ec0",
  1552 => x"fdc049eb",
  1553 => x"86c487d2",
  1554 => x"c5c187fe",
  1555 => x"1ec087c3",
  1556 => x"49f6e1c1",
  1557 => x"87c0fdc0",
  1558 => x"d4c11ec0",
  1559 => x"497087e8",
  1560 => x"87f4fcc0",
  1561 => x"f887c8c3",
  1562 => x"534f268e",
  1563 => x"61662044",
  1564 => x"64656c69",
  1565 => x"6f42002e",
  1566 => x"6e69746f",
  1567 => x"2e2e2e67",
  1568 => x"f1c01e00",
  1569 => x"87fa87fb",
  1570 => x"c31e4f26",
  1571 => x"c048ecc8",
  1572 => x"e8c8c378",
  1573 => x"fd78c048",
  1574 => x"87e587fc",
  1575 => x"4f2648c0",
  1576 => x"78452080",
  1577 => x"80007469",
  1578 => x"63614220",
  1579 => x"1264006b",
  1580 => x"32410000",
  1581 => x"00000000",
  1582 => x"00126400",
  1583 => x"00325f00",
  1584 => x"00000000",
  1585 => x"00001264",
  1586 => x"0000327d",
  1587 => x"64000000",
  1588 => x"9b000012",
  1589 => x"00000032",
  1590 => x"12640000",
  1591 => x"32b90000",
  1592 => x"00000000",
  1593 => x"00126400",
  1594 => x"0032d700",
  1595 => x"00000000",
  1596 => x"00001264",
  1597 => x"000032f5",
  1598 => x"64000000",
  1599 => x"00000012",
  1600 => x"00000000",
  1601 => x"12e80000",
  1602 => x"00000000",
  1603 => x"00000000",
  1604 => x"616f4c00",
  1605 => x"2e2a2064",
  1606 => x"f0fe1e00",
  1607 => x"cd78c048",
  1608 => x"26097909",
  1609 => x"fe1e1e4f",
  1610 => x"487ebff0",
  1611 => x"1e4f2626",
  1612 => x"c148f0fe",
  1613 => x"1e4f2678",
  1614 => x"c048f0fe",
  1615 => x"1e4f2678",
  1616 => x"52c04a71",
  1617 => x"0e4f2652",
  1618 => x"5d5c5b5e",
  1619 => x"7186f40e",
  1620 => x"7e6d974d",
  1621 => x"974ca5c1",
  1622 => x"a6c8486c",
  1623 => x"c4486e58",
  1624 => x"c505a866",
  1625 => x"c048ff87",
  1626 => x"caff87e6",
  1627 => x"49a5c287",
  1628 => x"714b6c97",
  1629 => x"6b974ba3",
  1630 => x"7e6c974b",
  1631 => x"80c1486e",
  1632 => x"c758a6c8",
  1633 => x"58a6cc98",
  1634 => x"fe7c9770",
  1635 => x"487387e1",
  1636 => x"4d268ef4",
  1637 => x"4b264c26",
  1638 => x"5e0e4f26",
  1639 => x"f40e5c5b",
  1640 => x"d84c7186",
  1641 => x"ffc34a66",
  1642 => x"4ba4c29a",
  1643 => x"73496c97",
  1644 => x"517249a1",
  1645 => x"6e7e6c97",
  1646 => x"c880c148",
  1647 => x"98c758a6",
  1648 => x"7058a6cc",
  1649 => x"ff8ef454",
  1650 => x"1e1e87ca",
  1651 => x"e087e8fd",
  1652 => x"c0494abf",
  1653 => x"0299c0e0",
  1654 => x"1e7287cb",
  1655 => x"49d3ccc3",
  1656 => x"c487f7fe",
  1657 => x"87fdfc86",
  1658 => x"c2fd7e70",
  1659 => x"4f262687",
  1660 => x"d3ccc31e",
  1661 => x"87c7fd49",
  1662 => x"49cae7c1",
  1663 => x"c587dafc",
  1664 => x"4f2687d0",
  1665 => x"5c5b5e0e",
  1666 => x"cdc30e5d",
  1667 => x"c14abfe6",
  1668 => x"49bfd8e9",
  1669 => x"71bc724c",
  1670 => x"87dbfc4d",
  1671 => x"49744bc0",
  1672 => x"d50299d0",
  1673 => x"d0497587",
  1674 => x"c01e7199",
  1675 => x"e1efc11e",
  1676 => x"1282734a",
  1677 => x"87e4c049",
  1678 => x"2cc186c8",
  1679 => x"abc8832d",
  1680 => x"87daff04",
  1681 => x"c187e8fb",
  1682 => x"c348d8e9",
  1683 => x"78bfe6cd",
  1684 => x"4c264d26",
  1685 => x"4f264b26",
  1686 => x"00000000",
  1687 => x"48d0ff1e",
  1688 => x"ff78e1c8",
  1689 => x"78c548d4",
  1690 => x"c30266c4",
  1691 => x"78e0c387",
  1692 => x"c60266c8",
  1693 => x"48d4ff87",
  1694 => x"ff78f0c3",
  1695 => x"787148d4",
  1696 => x"c848d0ff",
  1697 => x"e0c078e1",
  1698 => x"0e4f2678",
  1699 => x"0e5c5b5e",
  1700 => x"ccc34c71",
  1701 => x"eefa49d3",
  1702 => x"c04a7087",
  1703 => x"c204aab7",
  1704 => x"e0c387e3",
  1705 => x"87c905aa",
  1706 => x"48ceedc1",
  1707 => x"d4c278c1",
  1708 => x"aaf0c387",
  1709 => x"c187c905",
  1710 => x"c148caed",
  1711 => x"87f5c178",
  1712 => x"bfceedc1",
  1713 => x"7287c702",
  1714 => x"b3c0c24b",
  1715 => x"4b7287c2",
  1716 => x"d1059c74",
  1717 => x"caedc187",
  1718 => x"edc11ebf",
  1719 => x"721ebfce",
  1720 => x"87f8fd49",
  1721 => x"edc186c8",
  1722 => x"c002bfca",
  1723 => x"497387e0",
  1724 => x"9129b7c4",
  1725 => x"81e1eec1",
  1726 => x"9acf4a73",
  1727 => x"48c192c2",
  1728 => x"4a703072",
  1729 => x"4872baff",
  1730 => x"79709869",
  1731 => x"497387db",
  1732 => x"9129b7c4",
  1733 => x"81e1eec1",
  1734 => x"9acf4a73",
  1735 => x"48c392c2",
  1736 => x"4a703072",
  1737 => x"70b06948",
  1738 => x"ceedc179",
  1739 => x"c178c048",
  1740 => x"c048caed",
  1741 => x"d3ccc378",
  1742 => x"87cbf849",
  1743 => x"b7c04a70",
  1744 => x"ddfd03aa",
  1745 => x"fc48c087",
  1746 => x"000087c8",
  1747 => x"00000000",
  1748 => x"c01e0000",
  1749 => x"c449724a",
  1750 => x"e1eec191",
  1751 => x"c179c081",
  1752 => x"aab7d082",
  1753 => x"2687ee04",
  1754 => x"5b5e0e4f",
  1755 => x"710e5d5c",
  1756 => x"87c3f74d",
  1757 => x"b7c44a75",
  1758 => x"eec1922a",
  1759 => x"4c7582e1",
  1760 => x"94c29ccf",
  1761 => x"744b496a",
  1762 => x"c29bc32b",
  1763 => x"70307448",
  1764 => x"74bcff4c",
  1765 => x"70987148",
  1766 => x"87d3f67a",
  1767 => x"effa4873",
  1768 => x"00000087",
  1769 => x"00000000",
  1770 => x"00000000",
  1771 => x"00000000",
  1772 => x"00000000",
  1773 => x"00000000",
  1774 => x"00000000",
  1775 => x"00000000",
  1776 => x"00000000",
  1777 => x"00000000",
  1778 => x"00000000",
  1779 => x"00000000",
  1780 => x"00000000",
  1781 => x"00000000",
  1782 => x"00000000",
  1783 => x"00000000",
  1784 => x"261e1600",
  1785 => x"3d362e25",
  1786 => x"d0ff1e3e",
  1787 => x"78e1c848",
  1788 => x"d4ff4871",
  1789 => x"66c47808",
  1790 => x"08d4ff48",
  1791 => x"1e4f2678",
  1792 => x"66c44a71",
  1793 => x"49721e49",
  1794 => x"ff87deff",
  1795 => x"e0c048d0",
  1796 => x"4f262678",
  1797 => x"c24a711e",
  1798 => x"c303aab7",
  1799 => x"87c28287",
  1800 => x"66c482ce",
  1801 => x"ff49721e",
  1802 => x"262687d5",
  1803 => x"d4ff1e4f",
  1804 => x"7affc34a",
  1805 => x"c848d0ff",
  1806 => x"7ade78e1",
  1807 => x"bfddccc3",
  1808 => x"c848497a",
  1809 => x"717a7028",
  1810 => x"7028d048",
  1811 => x"d848717a",
  1812 => x"ff7a7028",
  1813 => x"e0c048d0",
  1814 => x"0e4f2678",
  1815 => x"5d5c5b5e",
  1816 => x"c34c710e",
  1817 => x"4dbfddcc",
  1818 => x"d02b744b",
  1819 => x"83c19b66",
  1820 => x"04ab66d4",
  1821 => x"4bc087c2",
  1822 => x"66d04a74",
  1823 => x"ff317249",
  1824 => x"739975b9",
  1825 => x"70307248",
  1826 => x"b071484a",
  1827 => x"58e1ccc3",
  1828 => x"2687dafe",
  1829 => x"264c264d",
  1830 => x"0e4f264b",
  1831 => x"5d5c5b5e",
  1832 => x"4c711e0e",
  1833 => x"4be1ccc3",
  1834 => x"f4c04ac0",
  1835 => x"d4d0fe49",
  1836 => x"c31e7487",
  1837 => x"fe49e1cc",
  1838 => x"c487ccee",
  1839 => x"02987086",
  1840 => x"c487eac0",
  1841 => x"1e4da61e",
  1842 => x"49e1ccc3",
  1843 => x"87fdf3fe",
  1844 => x"987086c8",
  1845 => x"7587d602",
  1846 => x"e3f4c14a",
  1847 => x"fe4bc449",
  1848 => x"7087c7ce",
  1849 => x"87ca0298",
  1850 => x"edc048c0",
  1851 => x"c048c087",
  1852 => x"f3c087e8",
  1853 => x"87c4c187",
  1854 => x"c8029870",
  1855 => x"87fcc087",
  1856 => x"f8059870",
  1857 => x"c1cdc387",
  1858 => x"87cc02bf",
  1859 => x"48ddccc3",
  1860 => x"bfc1cdc3",
  1861 => x"87d5fc78",
  1862 => x"262648c1",
  1863 => x"264c264d",
  1864 => x"5b4f264b",
  1865 => x"00435241",
  1866 => x"c31ec01e",
  1867 => x"fe49e1cc",
  1868 => x"c387f3f0",
  1869 => x"c048f9cc",
  1870 => x"4f262678",
  1871 => x"5c5b5e0e",
  1872 => x"86f40e5d",
  1873 => x"c048a6c4",
  1874 => x"f9ccc378",
  1875 => x"b7c348bf",
  1876 => x"87d103a8",
  1877 => x"bff9ccc3",
  1878 => x"c380c148",
  1879 => x"c058fdcc",
  1880 => x"e2c648fb",
  1881 => x"e1ccc387",
  1882 => x"f4f5fe49",
  1883 => x"c34c7087",
  1884 => x"4abff9cc",
  1885 => x"d8028ac3",
  1886 => x"028ac187",
  1887 => x"8a87cbc5",
  1888 => x"87f6c202",
  1889 => x"cdc1028a",
  1890 => x"c3028a87",
  1891 => x"e1c587e2",
  1892 => x"754dc087",
  1893 => x"c192c44a",
  1894 => x"c382e5fc",
  1895 => x"7548f5cc",
  1896 => x"6e7e7080",
  1897 => x"494bbf97",
  1898 => x"c1486e4b",
  1899 => x"816a50a3",
  1900 => x"a6cc4811",
  1901 => x"02ac7058",
  1902 => x"486e87c4",
  1903 => x"66c850c0",
  1904 => x"c387c705",
  1905 => x"c448f9cc",
  1906 => x"85c178a5",
  1907 => x"04adb7c4",
  1908 => x"c487c0ff",
  1909 => x"cdc387dc",
  1910 => x"c848bfc5",
  1911 => x"d101a8b7",
  1912 => x"02acca87",
  1913 => x"accd87cc",
  1914 => x"c087c702",
  1915 => x"c003acb7",
  1916 => x"cdc387f3",
  1917 => x"c84bbfc5",
  1918 => x"d203abb7",
  1919 => x"c9cdc387",
  1920 => x"c0817349",
  1921 => x"83c151e0",
  1922 => x"04abb7c8",
  1923 => x"c387eeff",
  1924 => x"c148d1cd",
  1925 => x"cfc150d2",
  1926 => x"50cdc150",
  1927 => x"80e450c0",
  1928 => x"cdc378c3",
  1929 => x"c5cdc387",
  1930 => x"c14849bf",
  1931 => x"c9cdc380",
  1932 => x"a0c44858",
  1933 => x"c2517481",
  1934 => x"f0c087f8",
  1935 => x"da04acb7",
  1936 => x"b7f9c087",
  1937 => x"87d301ac",
  1938 => x"bffdccc3",
  1939 => x"7491ca49",
  1940 => x"8af0c04a",
  1941 => x"48fdccc3",
  1942 => x"ca78a172",
  1943 => x"c6c002ac",
  1944 => x"05accd87",
  1945 => x"c387cbc2",
  1946 => x"c348f9cc",
  1947 => x"87c2c278",
  1948 => x"acb7f0c0",
  1949 => x"c087db04",
  1950 => x"01acb7f9",
  1951 => x"c387d3c0",
  1952 => x"49bfc1cd",
  1953 => x"4a7491d0",
  1954 => x"c38af0c0",
  1955 => x"7248c1cd",
  1956 => x"c1c178a1",
  1957 => x"c004acb7",
  1958 => x"c6c187db",
  1959 => x"c001acb7",
  1960 => x"cdc387d3",
  1961 => x"d049bfc1",
  1962 => x"c04a7491",
  1963 => x"cdc38af7",
  1964 => x"a17248c1",
  1965 => x"02acca78",
  1966 => x"cd87c6c0",
  1967 => x"f1c005ac",
  1968 => x"f9ccc387",
  1969 => x"c078c348",
  1970 => x"e2c087e8",
  1971 => x"c9c005ac",
  1972 => x"48a6c487",
  1973 => x"c078fbc0",
  1974 => x"acca87d8",
  1975 => x"87c6c002",
  1976 => x"c005accd",
  1977 => x"ccc387c9",
  1978 => x"78c348f9",
  1979 => x"c887c3c0",
  1980 => x"b7c05ca6",
  1981 => x"c4c003ac",
  1982 => x"cac04887",
  1983 => x"0266c487",
  1984 => x"4887c6f9",
  1985 => x"f499ffc3",
  1986 => x"87cff88e",
  1987 => x"464e4f43",
  1988 => x"4f4d003d",
  1989 => x"414e0044",
  1990 => x"4400454d",
  1991 => x"55414645",
  1992 => x"303d544c",
  1993 => x"001f0c00",
  1994 => x"001f1200",
  1995 => x"001f1600",
  1996 => x"001f1b00",
  1997 => x"d0ff1e00",
  1998 => x"78c9c848",
  1999 => x"d4ff4871",
  2000 => x"4f267808",
  2001 => x"494a711e",
  2002 => x"d0ff87eb",
  2003 => x"2678c848",
  2004 => x"1e731e4f",
  2005 => x"cdc34b71",
  2006 => x"c302bfe1",
  2007 => x"87ebc287",
  2008 => x"c848d0ff",
  2009 => x"497378c9",
  2010 => x"ffb1e0c0",
  2011 => x"787148d4",
  2012 => x"48d5cdc3",
  2013 => x"66c878c0",
  2014 => x"c387c502",
  2015 => x"87c249ff",
  2016 => x"cdc349c0",
  2017 => x"66cc59dd",
  2018 => x"c587c602",
  2019 => x"c44ad5d5",
  2020 => x"ffffcf87",
  2021 => x"e1cdc34a",
  2022 => x"e1cdc35a",
  2023 => x"c478c148",
  2024 => x"264d2687",
  2025 => x"264b264c",
  2026 => x"5b5e0e4f",
  2027 => x"710e5d5c",
  2028 => x"ddcdc34a",
  2029 => x"9a724cbf",
  2030 => x"4987cb02",
  2031 => x"fdc191c8",
  2032 => x"83714bc7",
  2033 => x"c1c287c4",
  2034 => x"4dc04bc7",
  2035 => x"99744913",
  2036 => x"bfd9cdc3",
  2037 => x"48d4ffb9",
  2038 => x"b7c17871",
  2039 => x"b7c8852c",
  2040 => x"87e804ad",
  2041 => x"bfd5cdc3",
  2042 => x"c380c848",
  2043 => x"fe58d9cd",
  2044 => x"731e87ef",
  2045 => x"134b711e",
  2046 => x"cb029a4a",
  2047 => x"fe497287",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
