
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom2 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"4a",x"13",x"87",x"e7"),
     1 => (x"87",x"f5",x"05",x"9a"),
     2 => (x"1e",x"87",x"da",x"fe"),
     3 => (x"bf",x"d5",x"cd",x"c3"),
     4 => (x"d5",x"cd",x"c3",x"49"),
     5 => (x"78",x"a1",x"c1",x"48"),
     6 => (x"a9",x"b7",x"c0",x"c4"),
     7 => (x"ff",x"87",x"db",x"03"),
     8 => (x"cd",x"c3",x"48",x"d4"),
     9 => (x"c3",x"78",x"bf",x"d9"),
    10 => (x"49",x"bf",x"d5",x"cd"),
    11 => (x"48",x"d5",x"cd",x"c3"),
    12 => (x"c4",x"78",x"a1",x"c1"),
    13 => (x"04",x"a9",x"b7",x"c0"),
    14 => (x"d0",x"ff",x"87",x"e5"),
    15 => (x"c3",x"78",x"c8",x"48"),
    16 => (x"c0",x"48",x"e1",x"cd"),
    17 => (x"00",x"4f",x"26",x"78"),
    18 => (x"00",x"00",x"00",x"00"),
    19 => (x"00",x"00",x"00",x"00"),
    20 => (x"5f",x"5f",x"00",x"00"),
    21 => (x"00",x"00",x"00",x"00"),
    22 => (x"03",x"00",x"03",x"03"),
    23 => (x"14",x"00",x"00",x"03"),
    24 => (x"7f",x"14",x"7f",x"7f"),
    25 => (x"00",x"00",x"14",x"7f"),
    26 => (x"6b",x"6b",x"2e",x"24"),
    27 => (x"4c",x"00",x"12",x"3a"),
    28 => (x"6c",x"18",x"36",x"6a"),
    29 => (x"30",x"00",x"32",x"56"),
    30 => (x"77",x"59",x"4f",x"7e"),
    31 => (x"00",x"40",x"68",x"3a"),
    32 => (x"03",x"07",x"04",x"00"),
    33 => (x"00",x"00",x"00",x"00"),
    34 => (x"63",x"3e",x"1c",x"00"),
    35 => (x"00",x"00",x"00",x"41"),
    36 => (x"3e",x"63",x"41",x"00"),
    37 => (x"08",x"00",x"00",x"1c"),
    38 => (x"1c",x"1c",x"3e",x"2a"),
    39 => (x"00",x"08",x"2a",x"3e"),
    40 => (x"3e",x"3e",x"08",x"08"),
    41 => (x"00",x"00",x"08",x"08"),
    42 => (x"60",x"e0",x"80",x"00"),
    43 => (x"00",x"00",x"00",x"00"),
    44 => (x"08",x"08",x"08",x"08"),
    45 => (x"00",x"00",x"08",x"08"),
    46 => (x"60",x"60",x"00",x"00"),
    47 => (x"40",x"00",x"00",x"00"),
    48 => (x"0c",x"18",x"30",x"60"),
    49 => (x"00",x"01",x"03",x"06"),
    50 => (x"4d",x"59",x"7f",x"3e"),
    51 => (x"00",x"00",x"3e",x"7f"),
    52 => (x"7f",x"7f",x"06",x"04"),
    53 => (x"00",x"00",x"00",x"00"),
    54 => (x"59",x"71",x"63",x"42"),
    55 => (x"00",x"00",x"46",x"4f"),
    56 => (x"49",x"49",x"63",x"22"),
    57 => (x"18",x"00",x"36",x"7f"),
    58 => (x"7f",x"13",x"16",x"1c"),
    59 => (x"00",x"00",x"10",x"7f"),
    60 => (x"45",x"45",x"67",x"27"),
    61 => (x"00",x"00",x"39",x"7d"),
    62 => (x"49",x"4b",x"7e",x"3c"),
    63 => (x"00",x"00",x"30",x"79"),
    64 => (x"79",x"71",x"01",x"01"),
    65 => (x"00",x"00",x"07",x"0f"),
    66 => (x"49",x"49",x"7f",x"36"),
    67 => (x"00",x"00",x"36",x"7f"),
    68 => (x"69",x"49",x"4f",x"06"),
    69 => (x"00",x"00",x"1e",x"3f"),
    70 => (x"66",x"66",x"00",x"00"),
    71 => (x"00",x"00",x"00",x"00"),
    72 => (x"66",x"e6",x"80",x"00"),
    73 => (x"00",x"00",x"00",x"00"),
    74 => (x"14",x"14",x"08",x"08"),
    75 => (x"00",x"00",x"22",x"22"),
    76 => (x"14",x"14",x"14",x"14"),
    77 => (x"00",x"00",x"14",x"14"),
    78 => (x"14",x"14",x"22",x"22"),
    79 => (x"00",x"00",x"08",x"08"),
    80 => (x"59",x"51",x"03",x"02"),
    81 => (x"3e",x"00",x"06",x"0f"),
    82 => (x"55",x"5d",x"41",x"7f"),
    83 => (x"00",x"00",x"1e",x"1f"),
    84 => (x"09",x"09",x"7f",x"7e"),
    85 => (x"00",x"00",x"7e",x"7f"),
    86 => (x"49",x"49",x"7f",x"7f"),
    87 => (x"00",x"00",x"36",x"7f"),
    88 => (x"41",x"63",x"3e",x"1c"),
    89 => (x"00",x"00",x"41",x"41"),
    90 => (x"63",x"41",x"7f",x"7f"),
    91 => (x"00",x"00",x"1c",x"3e"),
    92 => (x"49",x"49",x"7f",x"7f"),
    93 => (x"00",x"00",x"41",x"41"),
    94 => (x"09",x"09",x"7f",x"7f"),
    95 => (x"00",x"00",x"01",x"01"),
    96 => (x"49",x"41",x"7f",x"3e"),
    97 => (x"00",x"00",x"7a",x"7b"),
    98 => (x"08",x"08",x"7f",x"7f"),
    99 => (x"00",x"00",x"7f",x"7f"),
   100 => (x"7f",x"7f",x"41",x"00"),
   101 => (x"00",x"00",x"00",x"41"),
   102 => (x"40",x"40",x"60",x"20"),
   103 => (x"7f",x"00",x"3f",x"7f"),
   104 => (x"36",x"1c",x"08",x"7f"),
   105 => (x"00",x"00",x"41",x"63"),
   106 => (x"40",x"40",x"7f",x"7f"),
   107 => (x"7f",x"00",x"40",x"40"),
   108 => (x"06",x"0c",x"06",x"7f"),
   109 => (x"7f",x"00",x"7f",x"7f"),
   110 => (x"18",x"0c",x"06",x"7f"),
   111 => (x"00",x"00",x"7f",x"7f"),
   112 => (x"41",x"41",x"7f",x"3e"),
   113 => (x"00",x"00",x"3e",x"7f"),
   114 => (x"09",x"09",x"7f",x"7f"),
   115 => (x"3e",x"00",x"06",x"0f"),
   116 => (x"7f",x"61",x"41",x"7f"),
   117 => (x"00",x"00",x"40",x"7e"),
   118 => (x"19",x"09",x"7f",x"7f"),
   119 => (x"00",x"00",x"66",x"7f"),
   120 => (x"59",x"4d",x"6f",x"26"),
   121 => (x"00",x"00",x"32",x"7b"),
   122 => (x"7f",x"7f",x"01",x"01"),
   123 => (x"00",x"00",x"01",x"01"),
   124 => (x"40",x"40",x"7f",x"3f"),
   125 => (x"00",x"00",x"3f",x"7f"),
   126 => (x"70",x"70",x"3f",x"0f"),
   127 => (x"7f",x"00",x"0f",x"3f"),
   128 => (x"30",x"18",x"30",x"7f"),
   129 => (x"41",x"00",x"7f",x"7f"),
   130 => (x"1c",x"1c",x"36",x"63"),
   131 => (x"01",x"41",x"63",x"36"),
   132 => (x"7c",x"7c",x"06",x"03"),
   133 => (x"61",x"01",x"03",x"06"),
   134 => (x"47",x"4d",x"59",x"71"),
   135 => (x"00",x"00",x"41",x"43"),
   136 => (x"41",x"7f",x"7f",x"00"),
   137 => (x"01",x"00",x"00",x"41"),
   138 => (x"18",x"0c",x"06",x"03"),
   139 => (x"00",x"40",x"60",x"30"),
   140 => (x"7f",x"41",x"41",x"00"),
   141 => (x"08",x"00",x"00",x"7f"),
   142 => (x"06",x"03",x"06",x"0c"),
   143 => (x"80",x"00",x"08",x"0c"),
   144 => (x"80",x"80",x"80",x"80"),
   145 => (x"00",x"00",x"80",x"80"),
   146 => (x"07",x"03",x"00",x"00"),
   147 => (x"00",x"00",x"00",x"04"),
   148 => (x"54",x"54",x"74",x"20"),
   149 => (x"00",x"00",x"78",x"7c"),
   150 => (x"44",x"44",x"7f",x"7f"),
   151 => (x"00",x"00",x"38",x"7c"),
   152 => (x"44",x"44",x"7c",x"38"),
   153 => (x"00",x"00",x"00",x"44"),
   154 => (x"44",x"44",x"7c",x"38"),
   155 => (x"00",x"00",x"7f",x"7f"),
   156 => (x"54",x"54",x"7c",x"38"),
   157 => (x"00",x"00",x"18",x"5c"),
   158 => (x"05",x"7f",x"7e",x"04"),
   159 => (x"00",x"00",x"00",x"05"),
   160 => (x"a4",x"a4",x"bc",x"18"),
   161 => (x"00",x"00",x"7c",x"fc"),
   162 => (x"04",x"04",x"7f",x"7f"),
   163 => (x"00",x"00",x"78",x"7c"),
   164 => (x"7d",x"3d",x"00",x"00"),
   165 => (x"00",x"00",x"00",x"40"),
   166 => (x"fd",x"80",x"80",x"80"),
   167 => (x"00",x"00",x"00",x"7d"),
   168 => (x"38",x"10",x"7f",x"7f"),
   169 => (x"00",x"00",x"44",x"6c"),
   170 => (x"7f",x"3f",x"00",x"00"),
   171 => (x"7c",x"00",x"00",x"40"),
   172 => (x"0c",x"18",x"0c",x"7c"),
   173 => (x"00",x"00",x"78",x"7c"),
   174 => (x"04",x"04",x"7c",x"7c"),
   175 => (x"00",x"00",x"78",x"7c"),
   176 => (x"44",x"44",x"7c",x"38"),
   177 => (x"00",x"00",x"38",x"7c"),
   178 => (x"24",x"24",x"fc",x"fc"),
   179 => (x"00",x"00",x"18",x"3c"),
   180 => (x"24",x"24",x"3c",x"18"),
   181 => (x"00",x"00",x"fc",x"fc"),
   182 => (x"04",x"04",x"7c",x"7c"),
   183 => (x"00",x"00",x"08",x"0c"),
   184 => (x"54",x"54",x"5c",x"48"),
   185 => (x"00",x"00",x"20",x"74"),
   186 => (x"44",x"7f",x"3f",x"04"),
   187 => (x"00",x"00",x"00",x"44"),
   188 => (x"40",x"40",x"7c",x"3c"),
   189 => (x"00",x"00",x"7c",x"7c"),
   190 => (x"60",x"60",x"3c",x"1c"),
   191 => (x"3c",x"00",x"1c",x"3c"),
   192 => (x"60",x"30",x"60",x"7c"),
   193 => (x"44",x"00",x"3c",x"7c"),
   194 => (x"38",x"10",x"38",x"6c"),
   195 => (x"00",x"00",x"44",x"6c"),
   196 => (x"60",x"e0",x"bc",x"1c"),
   197 => (x"00",x"00",x"1c",x"3c"),
   198 => (x"5c",x"74",x"64",x"44"),
   199 => (x"00",x"00",x"44",x"4c"),
   200 => (x"77",x"3e",x"08",x"08"),
   201 => (x"00",x"00",x"41",x"41"),
   202 => (x"7f",x"7f",x"00",x"00"),
   203 => (x"00",x"00",x"00",x"00"),
   204 => (x"3e",x"77",x"41",x"41"),
   205 => (x"02",x"00",x"08",x"08"),
   206 => (x"02",x"03",x"01",x"01"),
   207 => (x"7f",x"00",x"01",x"02"),
   208 => (x"7f",x"7f",x"7f",x"7f"),
   209 => (x"08",x"00",x"7f",x"7f"),
   210 => (x"3e",x"1c",x"1c",x"08"),
   211 => (x"7f",x"7f",x"7f",x"3e"),
   212 => (x"1c",x"3e",x"3e",x"7f"),
   213 => (x"00",x"08",x"08",x"1c"),
   214 => (x"7c",x"7c",x"18",x"10"),
   215 => (x"00",x"00",x"10",x"18"),
   216 => (x"7c",x"7c",x"30",x"10"),
   217 => (x"10",x"00",x"10",x"30"),
   218 => (x"78",x"60",x"60",x"30"),
   219 => (x"42",x"00",x"06",x"1e"),
   220 => (x"3c",x"18",x"3c",x"66"),
   221 => (x"78",x"00",x"42",x"66"),
   222 => (x"c6",x"c2",x"6a",x"38"),
   223 => (x"60",x"00",x"38",x"6c"),
   224 => (x"00",x"60",x"00",x"00"),
   225 => (x"0e",x"00",x"60",x"00"),
   226 => (x"5d",x"5c",x"5b",x"5e"),
   227 => (x"4c",x"71",x"1e",x"0e"),
   228 => (x"bf",x"f2",x"cd",x"c3"),
   229 => (x"c0",x"4b",x"c0",x"4d"),
   230 => (x"02",x"ab",x"74",x"1e"),
   231 => (x"a6",x"c4",x"87",x"c7"),
   232 => (x"c5",x"78",x"c0",x"48"),
   233 => (x"48",x"a6",x"c4",x"87"),
   234 => (x"66",x"c4",x"78",x"c1"),
   235 => (x"ee",x"49",x"73",x"1e"),
   236 => (x"86",x"c8",x"87",x"df"),
   237 => (x"ef",x"49",x"e0",x"c0"),
   238 => (x"a5",x"c4",x"87",x"ef"),
   239 => (x"f0",x"49",x"6a",x"4a"),
   240 => (x"c6",x"f1",x"87",x"f0"),
   241 => (x"c1",x"85",x"cb",x"87"),
   242 => (x"ab",x"b7",x"c8",x"83"),
   243 => (x"87",x"c7",x"ff",x"04"),
   244 => (x"26",x"4d",x"26",x"26"),
   245 => (x"26",x"4b",x"26",x"4c"),
   246 => (x"4a",x"71",x"1e",x"4f"),
   247 => (x"5a",x"f6",x"cd",x"c3"),
   248 => (x"48",x"f6",x"cd",x"c3"),
   249 => (x"fe",x"49",x"78",x"c7"),
   250 => (x"4f",x"26",x"87",x"dd"),
   251 => (x"71",x"1e",x"73",x"1e"),
   252 => (x"aa",x"b7",x"c0",x"4a"),
   253 => (x"c2",x"87",x"d3",x"03"),
   254 => (x"05",x"bf",x"c2",x"e0"),
   255 => (x"4b",x"c1",x"87",x"c4"),
   256 => (x"4b",x"c0",x"87",x"c2"),
   257 => (x"5b",x"c6",x"e0",x"c2"),
   258 => (x"e0",x"c2",x"87",x"c4"),
   259 => (x"e0",x"c2",x"5a",x"c6"),
   260 => (x"c1",x"4a",x"bf",x"c2"),
   261 => (x"a2",x"c0",x"c1",x"9a"),
   262 => (x"87",x"e8",x"ec",x"49"),
   263 => (x"bf",x"ea",x"df",x"c2"),
   264 => (x"c2",x"e0",x"c2",x"49"),
   265 => (x"48",x"fc",x"b1",x"bf"),
   266 => (x"e8",x"fe",x"78",x"71"),
   267 => (x"4a",x"71",x"1e",x"87"),
   268 => (x"72",x"1e",x"66",x"c4"),
   269 => (x"db",x"df",x"ff",x"49"),
   270 => (x"4f",x"26",x"26",x"87"),
   271 => (x"c2",x"e0",x"c2",x"1e"),
   272 => (x"e2",x"c0",x"49",x"bf"),
   273 => (x"cd",x"c3",x"87",x"f0"),
   274 => (x"bf",x"e8",x"48",x"ea"),
   275 => (x"e6",x"cd",x"c3",x"78"),
   276 => (x"78",x"bf",x"ec",x"48"),
   277 => (x"bf",x"ea",x"cd",x"c3"),
   278 => (x"ff",x"c3",x"49",x"4a"),
   279 => (x"2a",x"b7",x"c8",x"99"),
   280 => (x"b0",x"71",x"48",x"72"),
   281 => (x"58",x"f2",x"cd",x"c3"),
   282 => (x"5e",x"0e",x"4f",x"26"),
   283 => (x"0e",x"5d",x"5c",x"5b"),
   284 => (x"c7",x"ff",x"4b",x"71"),
   285 => (x"e5",x"cd",x"c3",x"87"),
   286 => (x"73",x"50",x"c0",x"48"),
   287 => (x"e8",x"db",x"ff",x"49"),
   288 => (x"4c",x"49",x"70",x"87"),
   289 => (x"ee",x"cb",x"9c",x"c2"),
   290 => (x"87",x"fe",x"cd",x"49"),
   291 => (x"c3",x"4d",x"49",x"70"),
   292 => (x"bf",x"97",x"e5",x"cd"),
   293 => (x"87",x"e4",x"c1",x"05"),
   294 => (x"c3",x"49",x"66",x"d0"),
   295 => (x"99",x"bf",x"ee",x"cd"),
   296 => (x"d4",x"87",x"d7",x"05"),
   297 => (x"cd",x"c3",x"49",x"66"),
   298 => (x"05",x"99",x"bf",x"e6"),
   299 => (x"49",x"73",x"87",x"cc"),
   300 => (x"87",x"f5",x"da",x"ff"),
   301 => (x"c1",x"02",x"98",x"70"),
   302 => (x"4c",x"c1",x"87",x"c2"),
   303 => (x"75",x"87",x"fd",x"fd"),
   304 => (x"87",x"d2",x"cd",x"49"),
   305 => (x"c6",x"02",x"98",x"70"),
   306 => (x"e5",x"cd",x"c3",x"87"),
   307 => (x"c3",x"50",x"c1",x"48"),
   308 => (x"bf",x"97",x"e5",x"cd"),
   309 => (x"87",x"e4",x"c0",x"05"),
   310 => (x"bf",x"ee",x"cd",x"c3"),
   311 => (x"99",x"66",x"d0",x"49"),
   312 => (x"87",x"d6",x"ff",x"05"),
   313 => (x"bf",x"e6",x"cd",x"c3"),
   314 => (x"99",x"66",x"d4",x"49"),
   315 => (x"87",x"ca",x"ff",x"05"),
   316 => (x"d9",x"ff",x"49",x"73"),
   317 => (x"98",x"70",x"87",x"f3"),
   318 => (x"87",x"fe",x"fe",x"05"),
   319 => (x"d0",x"fb",x"48",x"74"),
   320 => (x"5b",x"5e",x"0e",x"87"),
   321 => (x"f8",x"0e",x"5d",x"5c"),
   322 => (x"4c",x"4d",x"c0",x"86"),
   323 => (x"c4",x"7e",x"bf",x"ec"),
   324 => (x"cd",x"c3",x"48",x"a6"),
   325 => (x"c0",x"78",x"bf",x"f2"),
   326 => (x"f7",x"c1",x"1e",x"1e"),
   327 => (x"87",x"ca",x"fd",x"49"),
   328 => (x"98",x"70",x"86",x"c8"),
   329 => (x"87",x"f3",x"c0",x"02"),
   330 => (x"bf",x"ea",x"df",x"c2"),
   331 => (x"c1",x"87",x"c4",x"05"),
   332 => (x"c0",x"87",x"c2",x"7e"),
   333 => (x"ea",x"df",x"c2",x"7e"),
   334 => (x"ca",x"78",x"6e",x"48"),
   335 => (x"66",x"c4",x"1e",x"fc"),
   336 => (x"c4",x"87",x"c9",x"02"),
   337 => (x"de",x"c2",x"48",x"a6"),
   338 => (x"87",x"c7",x"78",x"c1"),
   339 => (x"c2",x"48",x"a6",x"c4"),
   340 => (x"c4",x"78",x"cc",x"de"),
   341 => (x"ff",x"c8",x"49",x"66"),
   342 => (x"c1",x"86",x"c4",x"87"),
   343 => (x"c7",x"1e",x"c0",x"1e"),
   344 => (x"87",x"c6",x"fc",x"49"),
   345 => (x"98",x"70",x"86",x"c8"),
   346 => (x"ff",x"87",x"ce",x"02"),
   347 => (x"87",x"fc",x"f9",x"49"),
   348 => (x"ff",x"49",x"da",x"c1"),
   349 => (x"c1",x"87",x"f2",x"d7"),
   350 => (x"e5",x"cd",x"c3",x"4d"),
   351 => (x"c3",x"02",x"bf",x"97"),
   352 => (x"87",x"e4",x"cf",x"87"),
   353 => (x"bf",x"ea",x"cd",x"c3"),
   354 => (x"c2",x"e0",x"c2",x"4b"),
   355 => (x"e4",x"c1",x"05",x"bf"),
   356 => (x"ea",x"df",x"c2",x"87"),
   357 => (x"f1",x"c0",x"02",x"bf"),
   358 => (x"48",x"a6",x"c4",x"87"),
   359 => (x"78",x"c0",x"c0",x"c8"),
   360 => (x"7e",x"ee",x"df",x"c2"),
   361 => (x"49",x"bf",x"97",x"6e"),
   362 => (x"80",x"c1",x"48",x"6e"),
   363 => (x"ff",x"71",x"7e",x"70"),
   364 => (x"70",x"87",x"f6",x"d6"),
   365 => (x"87",x"c3",x"02",x"98"),
   366 => (x"c4",x"b3",x"66",x"c4"),
   367 => (x"b7",x"c1",x"48",x"66"),
   368 => (x"58",x"a6",x"c8",x"28"),
   369 => (x"ff",x"05",x"98",x"70"),
   370 => (x"fd",x"c3",x"87",x"da"),
   371 => (x"d8",x"d6",x"ff",x"49"),
   372 => (x"49",x"fa",x"c3",x"87"),
   373 => (x"87",x"d1",x"d6",x"ff"),
   374 => (x"ff",x"c3",x"49",x"73"),
   375 => (x"c0",x"1e",x"71",x"99"),
   376 => (x"87",x"c9",x"f9",x"49"),
   377 => (x"b7",x"c8",x"49",x"73"),
   378 => (x"c1",x"1e",x"71",x"29"),
   379 => (x"87",x"fd",x"f8",x"49"),
   380 => (x"c7",x"c6",x"86",x"c8"),
   381 => (x"ee",x"cd",x"c3",x"87"),
   382 => (x"02",x"9b",x"4b",x"bf"),
   383 => (x"df",x"c2",x"87",x"df"),
   384 => (x"c8",x"49",x"bf",x"fe"),
   385 => (x"98",x"70",x"87",x"d0"),
   386 => (x"87",x"c4",x"c0",x"05"),
   387 => (x"87",x"d3",x"4b",x"c0"),
   388 => (x"c7",x"49",x"e0",x"c2"),
   389 => (x"e0",x"c2",x"87",x"f4"),
   390 => (x"c6",x"c0",x"58",x"c2"),
   391 => (x"fe",x"df",x"c2",x"87"),
   392 => (x"73",x"78",x"c0",x"48"),
   393 => (x"05",x"99",x"c2",x"49"),
   394 => (x"c3",x"87",x"cf",x"c0"),
   395 => (x"d4",x"ff",x"49",x"eb"),
   396 => (x"49",x"70",x"87",x"f7"),
   397 => (x"c0",x"02",x"99",x"c2"),
   398 => (x"4c",x"fb",x"87",x"c2"),
   399 => (x"99",x"c1",x"49",x"73"),
   400 => (x"87",x"cf",x"c0",x"05"),
   401 => (x"ff",x"49",x"f4",x"c3"),
   402 => (x"70",x"87",x"de",x"d4"),
   403 => (x"02",x"99",x"c2",x"49"),
   404 => (x"fa",x"87",x"c2",x"c0"),
   405 => (x"c8",x"49",x"73",x"4c"),
   406 => (x"cf",x"c0",x"05",x"99"),
   407 => (x"49",x"f5",x"c3",x"87"),
   408 => (x"87",x"c5",x"d4",x"ff"),
   409 => (x"99",x"c2",x"49",x"70"),
   410 => (x"87",x"d6",x"c0",x"02"),
   411 => (x"bf",x"f6",x"cd",x"c3"),
   412 => (x"87",x"ca",x"c0",x"02"),
   413 => (x"c3",x"88",x"c1",x"48"),
   414 => (x"c0",x"58",x"fa",x"cd"),
   415 => (x"4c",x"ff",x"87",x"c2"),
   416 => (x"49",x"73",x"4d",x"c1"),
   417 => (x"c0",x"05",x"99",x"c4"),
   418 => (x"f2",x"c3",x"87",x"cf"),
   419 => (x"d8",x"d3",x"ff",x"49"),
   420 => (x"c2",x"49",x"70",x"87"),
   421 => (x"dc",x"c0",x"02",x"99"),
   422 => (x"f6",x"cd",x"c3",x"87"),
   423 => (x"c7",x"48",x"7e",x"bf"),
   424 => (x"c0",x"03",x"a8",x"b7"),
   425 => (x"48",x"6e",x"87",x"cb"),
   426 => (x"cd",x"c3",x"80",x"c1"),
   427 => (x"c2",x"c0",x"58",x"fa"),
   428 => (x"c1",x"4c",x"fe",x"87"),
   429 => (x"49",x"fd",x"c3",x"4d"),
   430 => (x"87",x"ed",x"d2",x"ff"),
   431 => (x"99",x"c2",x"49",x"70"),
   432 => (x"87",x"d5",x"c0",x"02"),
   433 => (x"bf",x"f6",x"cd",x"c3"),
   434 => (x"87",x"c9",x"c0",x"02"),
   435 => (x"48",x"f6",x"cd",x"c3"),
   436 => (x"c2",x"c0",x"78",x"c0"),
   437 => (x"c1",x"4c",x"fd",x"87"),
   438 => (x"49",x"fa",x"c3",x"4d"),
   439 => (x"87",x"c9",x"d2",x"ff"),
   440 => (x"99",x"c2",x"49",x"70"),
   441 => (x"87",x"d9",x"c0",x"02"),
   442 => (x"bf",x"f6",x"cd",x"c3"),
   443 => (x"a8",x"b7",x"c7",x"48"),
   444 => (x"87",x"c9",x"c0",x"03"),
   445 => (x"48",x"f6",x"cd",x"c3"),
   446 => (x"c2",x"c0",x"78",x"c7"),
   447 => (x"c1",x"4c",x"fc",x"87"),
   448 => (x"ac",x"b7",x"c0",x"4d"),
   449 => (x"87",x"d5",x"c0",x"03"),
   450 => (x"c1",x"48",x"66",x"c4"),
   451 => (x"7e",x"70",x"80",x"d8"),
   452 => (x"c0",x"02",x"bf",x"6e"),
   453 => (x"bf",x"6e",x"87",x"c7"),
   454 => (x"73",x"49",x"74",x"4b"),
   455 => (x"c3",x"1e",x"c0",x"0f"),
   456 => (x"da",x"c1",x"1e",x"f0"),
   457 => (x"87",x"c2",x"f5",x"49"),
   458 => (x"98",x"70",x"86",x"c8"),
   459 => (x"87",x"d9",x"c0",x"02"),
   460 => (x"bf",x"f6",x"cd",x"c3"),
   461 => (x"cb",x"49",x"6e",x"7e"),
   462 => (x"4a",x"66",x"c4",x"91"),
   463 => (x"02",x"6a",x"82",x"71"),
   464 => (x"6a",x"87",x"c6",x"c0"),
   465 => (x"73",x"49",x"6e",x"4b"),
   466 => (x"02",x"9d",x"75",x"0f"),
   467 => (x"c3",x"87",x"c8",x"c0"),
   468 => (x"49",x"bf",x"f6",x"cd"),
   469 => (x"c2",x"87",x"f0",x"f0"),
   470 => (x"02",x"bf",x"c6",x"e0"),
   471 => (x"49",x"87",x"dd",x"c0"),
   472 => (x"70",x"87",x"f3",x"c2"),
   473 => (x"d3",x"c0",x"02",x"98"),
   474 => (x"f6",x"cd",x"c3",x"87"),
   475 => (x"d6",x"f0",x"49",x"bf"),
   476 => (x"f1",x"49",x"c0",x"87"),
   477 => (x"e0",x"c2",x"87",x"f6"),
   478 => (x"78",x"c0",x"48",x"c6"),
   479 => (x"d0",x"f1",x"8e",x"f8"),
   480 => (x"79",x"6f",x"4a",x"87"),
   481 => (x"73",x"79",x"65",x"6b"),
   482 => (x"00",x"6e",x"6f",x"20"),
   483 => (x"6b",x"79",x"6f",x"4a"),
   484 => (x"20",x"73",x"79",x"65"),
   485 => (x"00",x"66",x"66",x"6f"),
   486 => (x"5c",x"5b",x"5e",x"0e"),
   487 => (x"71",x"1e",x"0e",x"5d"),
   488 => (x"f2",x"cd",x"c3",x"4c"),
   489 => (x"cd",x"c1",x"49",x"bf"),
   490 => (x"d1",x"c1",x"4d",x"a1"),
   491 => (x"74",x"7e",x"69",x"81"),
   492 => (x"87",x"cf",x"02",x"9c"),
   493 => (x"74",x"4b",x"a5",x"c4"),
   494 => (x"f2",x"cd",x"c3",x"7b"),
   495 => (x"d8",x"f0",x"49",x"bf"),
   496 => (x"74",x"7b",x"6e",x"87"),
   497 => (x"87",x"c4",x"05",x"9c"),
   498 => (x"87",x"c2",x"4b",x"c0"),
   499 => (x"49",x"73",x"4b",x"c1"),
   500 => (x"d4",x"87",x"d9",x"f0"),
   501 => (x"87",x"c8",x"02",x"66"),
   502 => (x"87",x"ee",x"c0",x"49"),
   503 => (x"87",x"c2",x"4a",x"70"),
   504 => (x"e0",x"c2",x"4a",x"c0"),
   505 => (x"ef",x"26",x"5a",x"ca"),
   506 => (x"00",x"00",x"87",x"e7"),
   507 => (x"12",x"58",x"00",x"00"),
   508 => (x"1b",x"1d",x"14",x"11"),
   509 => (x"59",x"5a",x"23",x"1c"),
   510 => (x"f2",x"f5",x"94",x"91"),
   511 => (x"00",x"00",x"f4",x"eb"),
   512 => (x"00",x"00",x"00",x"00"),
   513 => (x"00",x"00",x"00",x"00"),
   514 => (x"71",x"1e",x"00",x"00"),
   515 => (x"bf",x"c8",x"ff",x"4a"),
   516 => (x"48",x"a1",x"72",x"49"),
   517 => (x"ff",x"1e",x"4f",x"26"),
   518 => (x"fe",x"89",x"bf",x"c8"),
   519 => (x"c0",x"c0",x"c0",x"c0"),
   520 => (x"c4",x"01",x"a9",x"c0"),
   521 => (x"c2",x"4a",x"c0",x"87"),
   522 => (x"72",x"4a",x"c1",x"87"),
   523 => (x"0e",x"4f",x"26",x"48"),
   524 => (x"5d",x"5c",x"5b",x"5e"),
   525 => (x"4d",x"71",x"1e",x"0e"),
   526 => (x"75",x"4b",x"d4",x"ff"),
   527 => (x"fa",x"cd",x"c3",x"1e"),
   528 => (x"c2",x"c0",x"fe",x"49"),
   529 => (x"70",x"86",x"c4",x"87"),
   530 => (x"c3",x"02",x"6e",x"7e"),
   531 => (x"ce",x"c3",x"87",x"ff"),
   532 => (x"75",x"4c",x"bf",x"c2"),
   533 => (x"f0",x"d9",x"fe",x"49"),
   534 => (x"05",x"a8",x"de",x"87"),
   535 => (x"75",x"87",x"eb",x"c0"),
   536 => (x"f6",x"d0",x"ff",x"49"),
   537 => (x"02",x"98",x"70",x"87"),
   538 => (x"cc",x"c3",x"87",x"db"),
   539 => (x"c0",x"1e",x"bf",x"fd"),
   540 => (x"ce",x"ff",x"49",x"e1"),
   541 => (x"86",x"c4",x"87",x"c9"),
   542 => (x"48",x"e7",x"e5",x"c2"),
   543 => (x"cd",x"c3",x"50",x"c0"),
   544 => (x"ea",x"fe",x"49",x"c9"),
   545 => (x"c3",x"48",x"c1",x"87"),
   546 => (x"d0",x"ff",x"87",x"c5"),
   547 => (x"78",x"c5",x"c8",x"48"),
   548 => (x"c0",x"7b",x"d6",x"c1"),
   549 => (x"bf",x"97",x"6e",x"4a"),
   550 => (x"c1",x"48",x"6e",x"7b"),
   551 => (x"c1",x"7e",x"70",x"80"),
   552 => (x"b7",x"e0",x"c0",x"82"),
   553 => (x"ec",x"ff",x"04",x"aa"),
   554 => (x"48",x"d0",x"ff",x"87"),
   555 => (x"c5",x"c8",x"78",x"c4"),
   556 => (x"7b",x"d3",x"c1",x"78"),
   557 => (x"78",x"c4",x"7b",x"c1"),
   558 => (x"c1",x"02",x"9c",x"74"),
   559 => (x"fb",x"c2",x"87",x"fd"),
   560 => (x"c0",x"c8",x"7e",x"f6"),
   561 => (x"b7",x"c0",x"8c",x"4d"),
   562 => (x"87",x"c6",x"03",x"ac"),
   563 => (x"4d",x"a4",x"c0",x"c8"),
   564 => (x"c8",x"c3",x"4c",x"c0"),
   565 => (x"49",x"bf",x"97",x"e7"),
   566 => (x"d2",x"02",x"99",x"d0"),
   567 => (x"c3",x"1e",x"c0",x"87"),
   568 => (x"fe",x"49",x"fa",x"cd"),
   569 => (x"c4",x"87",x"fc",x"c0"),
   570 => (x"4a",x"49",x"70",x"86"),
   571 => (x"c2",x"87",x"ef",x"c0"),
   572 => (x"c3",x"1e",x"f6",x"fb"),
   573 => (x"fe",x"49",x"fa",x"cd"),
   574 => (x"c4",x"87",x"e8",x"c0"),
   575 => (x"4a",x"49",x"70",x"86"),
   576 => (x"c8",x"48",x"d0",x"ff"),
   577 => (x"d4",x"c1",x"78",x"c5"),
   578 => (x"bf",x"97",x"6e",x"7b"),
   579 => (x"c1",x"48",x"6e",x"7b"),
   580 => (x"c1",x"7e",x"70",x"80"),
   581 => (x"f0",x"ff",x"05",x"8d"),
   582 => (x"48",x"d0",x"ff",x"87"),
   583 => (x"9a",x"72",x"78",x"c4"),
   584 => (x"87",x"c5",x"c0",x"05"),
   585 => (x"e6",x"c0",x"48",x"c0"),
   586 => (x"c3",x"1e",x"c1",x"87"),
   587 => (x"fd",x"49",x"fa",x"cd"),
   588 => (x"c4",x"87",x"cf",x"fe"),
   589 => (x"05",x"9c",x"74",x"86"),
   590 => (x"ff",x"87",x"c3",x"fe"),
   591 => (x"c5",x"c8",x"48",x"d0"),
   592 => (x"7b",x"d3",x"c1",x"78"),
   593 => (x"78",x"c4",x"7b",x"c0"),
   594 => (x"c2",x"c0",x"48",x"c1"),
   595 => (x"26",x"48",x"c0",x"87"),
   596 => (x"4c",x"26",x"4d",x"26"),
   597 => (x"4f",x"26",x"4b",x"26"),
   598 => (x"c4",x"4a",x"71",x"1e"),
   599 => (x"87",x"c5",x"05",x"66"),
   600 => (x"ca",x"fb",x"49",x"72"),
   601 => (x"00",x"4f",x"26",x"87"),
   602 => (x"f6",x"e6",x"c2",x"1e"),
   603 => (x"b9",x"c1",x"49",x"bf"),
   604 => (x"59",x"fa",x"e6",x"c2"),
   605 => (x"c3",x"48",x"d4",x"ff"),
   606 => (x"d0",x"ff",x"78",x"ff"),
   607 => (x"78",x"e1",x"c8",x"48"),
   608 => (x"c1",x"48",x"d4",x"ff"),
   609 => (x"71",x"31",x"c4",x"78"),
   610 => (x"48",x"d0",x"ff",x"78"),
   611 => (x"26",x"78",x"e0",x"c0"),
   612 => (x"e6",x"c2",x"1e",x"4f"),
   613 => (x"cd",x"c3",x"1e",x"ea"),
   614 => (x"fa",x"fd",x"49",x"fa"),
   615 => (x"86",x"c4",x"87",x"e9"),
   616 => (x"c3",x"02",x"98",x"70"),
   617 => (x"87",x"c0",x"ff",x"87"),
   618 => (x"35",x"31",x"4f",x"26"),
   619 => (x"20",x"5a",x"48",x"4b"),
   620 => (x"46",x"43",x"20",x"20"),
   621 => (x"00",x"00",x"00",x"47"),
   622 => (x"fe",x"1e",x"00",x"00"),
   623 => (x"c4",x"87",x"f8",x"fd"),
   624 => (x"c0",x"c2",x"49",x"66"),
   625 => (x"87",x"cd",x"02",x"99"),
   626 => (x"c3",x"1e",x"e0",x"c3"),
   627 => (x"fe",x"49",x"d3",x"cc"),
   628 => (x"c4",x"87",x"c7",x"ff"),
   629 => (x"49",x"66",x"c4",x"86"),
   630 => (x"02",x"99",x"c0",x"c4"),
   631 => (x"f0",x"c3",x"87",x"cd"),
   632 => (x"d3",x"cc",x"c3",x"1e"),
   633 => (x"f1",x"fe",x"fe",x"49"),
   634 => (x"c4",x"86",x"c4",x"87"),
   635 => (x"ff",x"c1",x"49",x"66"),
   636 => (x"c3",x"1e",x"71",x"99"),
   637 => (x"fe",x"49",x"d3",x"cc"),
   638 => (x"fe",x"87",x"df",x"fe"),
   639 => (x"26",x"87",x"f0",x"fc"),
   640 => (x"5e",x"0e",x"4f",x"26"),
   641 => (x"0e",x"5d",x"5c",x"5b"),
   642 => (x"c0",x"86",x"d8",x"ff"),
   643 => (x"d2",x"ce",x"c3",x"7e"),
   644 => (x"81",x"c2",x"49",x"bf"),
   645 => (x"1e",x"72",x"1e",x"71"),
   646 => (x"db",x"fd",x"4a",x"c6"),
   647 => (x"48",x"71",x"87",x"e8"),
   648 => (x"49",x"26",x"4a",x"26"),
   649 => (x"c3",x"58",x"a6",x"c8"),
   650 => (x"49",x"bf",x"d2",x"ce"),
   651 => (x"1e",x"71",x"81",x"c4"),
   652 => (x"4a",x"c6",x"1e",x"72"),
   653 => (x"87",x"ce",x"db",x"fd"),
   654 => (x"4a",x"26",x"48",x"71"),
   655 => (x"a6",x"cc",x"49",x"26"),
   656 => (x"d3",x"f3",x"c2",x"58"),
   657 => (x"cd",x"f7",x"49",x"bf"),
   658 => (x"02",x"98",x"70",x"87"),
   659 => (x"c0",x"87",x"f9",x"c9"),
   660 => (x"f5",x"f6",x"49",x"e0"),
   661 => (x"c2",x"49",x"70",x"87"),
   662 => (x"c0",x"59",x"d7",x"f3"),
   663 => (x"c4",x"49",x"74",x"4c"),
   664 => (x"81",x"d0",x"fe",x"91"),
   665 => (x"49",x"74",x"4a",x"69"),
   666 => (x"bf",x"d2",x"ce",x"c3"),
   667 => (x"c3",x"91",x"c4",x"81"),
   668 => (x"72",x"81",x"de",x"ce"),
   669 => (x"d2",x"02",x"9a",x"79"),
   670 => (x"c1",x"49",x"72",x"87"),
   671 => (x"6e",x"9a",x"71",x"89"),
   672 => (x"70",x"80",x"c1",x"48"),
   673 => (x"05",x"9a",x"72",x"7e"),
   674 => (x"c1",x"87",x"ee",x"ff"),
   675 => (x"ac",x"b7",x"c2",x"84"),
   676 => (x"87",x"c9",x"ff",x"04"),
   677 => (x"fc",x"c0",x"48",x"6e"),
   678 => (x"c8",x"04",x"a8",x"b7"),
   679 => (x"4c",x"c0",x"87",x"ea"),
   680 => (x"66",x"c4",x"4a",x"74"),
   681 => (x"c3",x"92",x"c4",x"82"),
   682 => (x"74",x"82",x"de",x"ce"),
   683 => (x"81",x"66",x"c8",x"49"),
   684 => (x"ce",x"c3",x"91",x"c4"),
   685 => (x"4a",x"6a",x"81",x"de"),
   686 => (x"b9",x"72",x"49",x"69"),
   687 => (x"ce",x"c3",x"4b",x"74"),
   688 => (x"c4",x"83",x"bf",x"d2"),
   689 => (x"de",x"ce",x"c3",x"93"),
   690 => (x"72",x"ba",x"6b",x"83"),
   691 => (x"d4",x"98",x"71",x"48"),
   692 => (x"49",x"74",x"58",x"a6"),
   693 => (x"bf",x"d2",x"ce",x"c3"),
   694 => (x"c3",x"91",x"c4",x"81"),
   695 => (x"69",x"81",x"de",x"ce"),
   696 => (x"48",x"a6",x"d4",x"7e"),
   697 => (x"a6",x"d0",x"78",x"c0"),
   698 => (x"4c",x"ff",x"c3",x"5c"),
   699 => (x"df",x"49",x"66",x"d0"),
   700 => (x"e2",x"c6",x"02",x"29"),
   701 => (x"4a",x"66",x"cc",x"87"),
   702 => (x"d4",x"92",x"e0",x"c0"),
   703 => (x"ff",x"c0",x"82",x"66"),
   704 => (x"70",x"88",x"72",x"48"),
   705 => (x"48",x"a6",x"d8",x"4a"),
   706 => (x"80",x"c4",x"78",x"c0"),
   707 => (x"49",x"6e",x"78",x"c0"),
   708 => (x"e4",x"c0",x"29",x"df"),
   709 => (x"ce",x"c3",x"59",x"a6"),
   710 => (x"78",x"c1",x"48",x"ce"),
   711 => (x"31",x"c3",x"49",x"72"),
   712 => (x"b1",x"72",x"2a",x"b7"),
   713 => (x"c4",x"99",x"ff",x"c0"),
   714 => (x"ce",x"f7",x"c2",x"91"),
   715 => (x"6d",x"85",x"71",x"4d"),
   716 => (x"c0",x"c4",x"49",x"4b"),
   717 => (x"d7",x"02",x"99",x"c0"),
   718 => (x"66",x"e0",x"c0",x"87"),
   719 => (x"87",x"c7",x"c0",x"02"),
   720 => (x"78",x"c0",x"80",x"c8"),
   721 => (x"c3",x"87",x"d0",x"c5"),
   722 => (x"c1",x"48",x"d6",x"ce"),
   723 => (x"87",x"c7",x"c5",x"78"),
   724 => (x"02",x"66",x"e0",x"c0"),
   725 => (x"49",x"73",x"87",x"d8"),
   726 => (x"99",x"c0",x"c0",x"c2"),
   727 => (x"87",x"c3",x"c0",x"02"),
   728 => (x"6d",x"2b",x"b7",x"d0"),
   729 => (x"ff",x"ff",x"fd",x"48"),
   730 => (x"c0",x"7d",x"70",x"98"),
   731 => (x"ce",x"c3",x"87",x"fa"),
   732 => (x"c0",x"02",x"bf",x"d6"),
   733 => (x"48",x"73",x"87",x"f2"),
   734 => (x"c0",x"28",x"b7",x"d0"),
   735 => (x"70",x"58",x"a6",x"e8"),
   736 => (x"e3",x"c0",x"02",x"98"),
   737 => (x"da",x"ce",x"c3",x"87"),
   738 => (x"e0",x"c0",x"49",x"bf"),
   739 => (x"c0",x"02",x"99",x"c0"),
   740 => (x"49",x"70",x"87",x"ca"),
   741 => (x"99",x"c0",x"e0",x"c0"),
   742 => (x"87",x"cc",x"c0",x"02"),
   743 => (x"c0",x"c2",x"48",x"6d"),
   744 => (x"7d",x"70",x"b0",x"c0"),
   745 => (x"4b",x"66",x"e4",x"c0"),
   746 => (x"c0",x"c8",x"49",x"73"),
   747 => (x"c2",x"02",x"99",x"c0"),
   748 => (x"ce",x"c3",x"87",x"c5"),
   749 => (x"cc",x"4a",x"bf",x"da"),
   750 => (x"c0",x"02",x"9a",x"c0"),
   751 => (x"c0",x"c4",x"87",x"cf"),
   752 => (x"d7",x"c0",x"02",x"8a"),
   753 => (x"c0",x"02",x"8a",x"87"),
   754 => (x"dc",x"c1",x"87",x"f8"),
   755 => (x"74",x"49",x"73",x"87"),
   756 => (x"c2",x"91",x"c2",x"99"),
   757 => (x"11",x"81",x"c2",x"f7"),
   758 => (x"87",x"db",x"c1",x"4b"),
   759 => (x"99",x"74",x"49",x"73"),
   760 => (x"f7",x"c2",x"91",x"c2"),
   761 => (x"81",x"c1",x"81",x"c2"),
   762 => (x"e0",x"c0",x"4b",x"11"),
   763 => (x"c8",x"c0",x"02",x"66"),
   764 => (x"48",x"a6",x"dc",x"87"),
   765 => (x"fe",x"c0",x"78",x"d2"),
   766 => (x"48",x"a6",x"d8",x"87"),
   767 => (x"c0",x"78",x"d2",x"c4"),
   768 => (x"49",x"73",x"87",x"f5"),
   769 => (x"91",x"c2",x"99",x"74"),
   770 => (x"81",x"c2",x"f7",x"c2"),
   771 => (x"4b",x"11",x"81",x"c1"),
   772 => (x"02",x"66",x"e0",x"c0"),
   773 => (x"dc",x"87",x"c9",x"c0"),
   774 => (x"d9",x"c1",x"48",x"a6"),
   775 => (x"87",x"d7",x"c0",x"78"),
   776 => (x"c5",x"48",x"a6",x"d8"),
   777 => (x"ce",x"c0",x"78",x"d9"),
   778 => (x"74",x"49",x"73",x"87"),
   779 => (x"c2",x"91",x"c2",x"99"),
   780 => (x"c1",x"81",x"c2",x"f7"),
   781 => (x"c0",x"4b",x"11",x"81"),
   782 => (x"c0",x"02",x"66",x"e0"),
   783 => (x"49",x"73",x"87",x"db"),
   784 => (x"fc",x"c7",x"b9",x"ff"),
   785 => (x"48",x"71",x"99",x"c0"),
   786 => (x"bf",x"da",x"ce",x"c3"),
   787 => (x"de",x"ce",x"c3",x"98"),
   788 => (x"c4",x"9b",x"74",x"58"),
   789 => (x"d3",x"c0",x"b3",x"c0"),
   790 => (x"c7",x"49",x"73",x"87"),
   791 => (x"71",x"99",x"c0",x"fc"),
   792 => (x"da",x"ce",x"c3",x"48"),
   793 => (x"ce",x"c3",x"b0",x"bf"),
   794 => (x"9b",x"74",x"58",x"de"),
   795 => (x"c0",x"02",x"66",x"d8"),
   796 => (x"c3",x"1e",x"87",x"ca"),
   797 => (x"f5",x"49",x"ce",x"ce"),
   798 => (x"86",x"c4",x"87",x"c0"),
   799 => (x"ce",x"c3",x"1e",x"73"),
   800 => (x"f5",x"f4",x"49",x"ce"),
   801 => (x"dc",x"86",x"c4",x"87"),
   802 => (x"ca",x"c0",x"02",x"66"),
   803 => (x"ce",x"c3",x"1e",x"87"),
   804 => (x"e5",x"f4",x"49",x"ce"),
   805 => (x"d0",x"86",x"c4",x"87"),
   806 => (x"30",x"c1",x"48",x"66"),
   807 => (x"6e",x"58",x"a6",x"d4"),
   808 => (x"70",x"30",x"c1",x"48"),
   809 => (x"48",x"66",x"d4",x"7e"),
   810 => (x"a6",x"d8",x"80",x"c1"),
   811 => (x"b7",x"e0",x"c0",x"58"),
   812 => (x"f7",x"f8",x"04",x"a8"),
   813 => (x"4c",x"66",x"cc",x"87"),
   814 => (x"b7",x"c2",x"84",x"c1"),
   815 => (x"df",x"f7",x"04",x"ac"),
   816 => (x"d2",x"ce",x"c3",x"87"),
   817 => (x"78",x"66",x"c4",x"48"),
   818 => (x"26",x"8e",x"d8",x"ff"),
   819 => (x"26",x"4c",x"26",x"4d"),
   820 => (x"00",x"4f",x"26",x"4b"),
   821 => (x"1e",x"00",x"00",x"00"),
   822 => (x"49",x"72",x"4a",x"c0"),
   823 => (x"ce",x"c3",x"91",x"c4"),
   824 => (x"79",x"ff",x"81",x"de"),
   825 => (x"b7",x"c6",x"82",x"c1"),
   826 => (x"87",x"ee",x"04",x"aa"),
   827 => (x"48",x"d2",x"ce",x"c3"),
   828 => (x"78",x"40",x"40",x"c0"),
   829 => (x"73",x"1e",x"4f",x"26"),
   830 => (x"f4",x"4b",x"71",x"1e"),
   831 => (x"49",x"73",x"87",x"c4"),
   832 => (x"87",x"c7",x"f6",x"fe"),
   833 => (x"0e",x"87",x"c8",x"ff"),
   834 => (x"0e",x"5c",x"5b",x"5e"),
   835 => (x"ff",x"4c",x"d4",x"ff"),
   836 => (x"c5",x"c8",x"4b",x"d0"),
   837 => (x"7c",x"d5",x"c1",x"7b"),
   838 => (x"c4",x"7c",x"66",x"cc"),
   839 => (x"7b",x"c5",x"c8",x"7b"),
   840 => (x"c1",x"7c",x"d3",x"c1"),
   841 => (x"c8",x"7b",x"c4",x"7c"),
   842 => (x"d4",x"c1",x"7b",x"c5"),
   843 => (x"b7",x"4a",x"c0",x"7c"),
   844 => (x"87",x"cb",x"06",x"a9"),
   845 => (x"c1",x"7c",x"ff",x"c3"),
   846 => (x"aa",x"b7",x"71",x"82"),
   847 => (x"c4",x"87",x"f5",x"04"),
   848 => (x"7b",x"c5",x"c8",x"7b"),
   849 => (x"c0",x"7c",x"d3",x"c1"),
   850 => (x"fd",x"7b",x"c4",x"7c"),
   851 => (x"73",x"1e",x"87",x"ff"),
   852 => (x"49",x"4b",x"71",x"1e"),
   853 => (x"e2",x"c1",x"91",x"cb"),
   854 => (x"82",x"71",x"4a",x"ee"),
   855 => (x"97",x"e5",x"cd",x"c3"),
   856 => (x"87",x"d3",x"02",x"bf"),
   857 => (x"11",x"49",x"a2",x"ca"),
   858 => (x"c1",x"87",x"cc",x"05"),
   859 => (x"49",x"c0",x"c8",x"1e"),
   860 => (x"c4",x"87",x"d4",x"fe"),
   861 => (x"73",x"87",x"cc",x"86"),
   862 => (x"f7",x"d4",x"fe",x"49"),
   863 => (x"fe",x"49",x"73",x"87"),
   864 => (x"fd",x"87",x"f1",x"d4"),
   865 => (x"73",x"1e",x"87",x"c9"),
   866 => (x"c2",x"4b",x"c0",x"1e"),
   867 => (x"ea",x"49",x"e3",x"f6"),
   868 => (x"98",x"70",x"87",x"dd"),
   869 => (x"c2",x"87",x"c4",x"05"),
   870 => (x"fc",x"4b",x"ef",x"f6"),
   871 => (x"48",x"73",x"87",x"f9"),
   872 => (x"53",x"87",x"ec",x"fc"),
   873 => (x"32",x"33",x"49",x"56"),
   874 => (x"52",x"20",x"20",x"38"),
   875 => (x"52",x"00",x"4d",x"4f"),
   876 => (x"6c",x"20",x"4d",x"4f"),
   877 => (x"69",x"64",x"61",x"6f"),
   878 => (x"66",x"20",x"67",x"6e"),
   879 => (x"65",x"6c",x"69",x"61"),
   880 => (x"eb",x"f4",x"00",x"64"),
   881 => (x"06",x"05",x"f5",x"f2"),
   882 => (x"0b",x"03",x"0c",x"04"),
   883 => (x"00",x"66",x"0a",x"83"),
   884 => (x"00",x"5a",x"00",x"fc"),
   885 => (x"80",x"00",x"00",x"da"),
   886 => (x"80",x"05",x"08",x"94"),
   887 => (x"80",x"02",x"00",x"78"),
   888 => (x"80",x"03",x"00",x"01"),
   889 => (x"80",x"04",x"00",x"09"),
   890 => (x"80",x"01",x"00",x"00"),
   891 => (x"00",x"26",x"08",x"91"),
   892 => (x"00",x"1d",x"00",x"04"),
   893 => (x"00",x"1c",x"00",x"00"),
   894 => (x"00",x"25",x"00",x"00"),
   895 => (x"00",x"1a",x"00",x"0c"),
   896 => (x"00",x"1b",x"00",x"00"),
   897 => (x"00",x"24",x"00",x"00"),
   898 => (x"01",x"12",x"00",x"00"),
   899 => (x"00",x"2e",x"00",x"00"),
   900 => (x"00",x"2d",x"00",x"03"),
   901 => (x"00",x"23",x"00",x"00"),
   902 => (x"00",x"36",x"00",x"00"),
   903 => (x"00",x"21",x"00",x"0b"),
   904 => (x"00",x"2b",x"00",x"00"),
   905 => (x"00",x"2c",x"00",x"00"),
   906 => (x"00",x"22",x"00",x"00"),
   907 => (x"00",x"3d",x"00",x"00"),
   908 => (x"00",x"35",x"00",x"6c"),
   909 => (x"00",x"34",x"00",x"00"),
   910 => (x"00",x"3e",x"00",x"00"),
   911 => (x"00",x"32",x"00",x"75"),
   912 => (x"00",x"33",x"00",x"00"),
   913 => (x"00",x"3c",x"00",x"00"),
   914 => (x"00",x"2a",x"00",x"6b"),
   915 => (x"00",x"46",x"00",x"00"),
   916 => (x"00",x"43",x"00",x"01"),
   917 => (x"00",x"3b",x"00",x"73"),
   918 => (x"00",x"45",x"00",x"69"),
   919 => (x"00",x"3a",x"00",x"09"),
   920 => (x"00",x"42",x"00",x"70"),
   921 => (x"00",x"44",x"00",x"72"),
   922 => (x"00",x"31",x"00",x"74"),
   923 => (x"00",x"55",x"00",x"00"),
   924 => (x"00",x"4d",x"00",x"00"),
   925 => (x"00",x"4b",x"00",x"7c"),
   926 => (x"00",x"7b",x"00",x"7a"),
   927 => (x"00",x"49",x"00",x"00"),
   928 => (x"00",x"4c",x"00",x"71"),
   929 => (x"00",x"54",x"00",x"84"),
   930 => (x"00",x"41",x"00",x"77"),
   931 => (x"00",x"61",x"00",x"00"),
   932 => (x"00",x"5b",x"00",x"00"),
   933 => (x"00",x"52",x"00",x"7c"),
   934 => (x"00",x"f1",x"00",x"00"),
   935 => (x"02",x"59",x"00",x"00"),
   936 => (x"00",x"0e",x"00",x"00"),
   937 => (x"00",x"5d",x"00",x"5d"),
   938 => (x"00",x"4a",x"00",x"00"),
   939 => (x"00",x"16",x"00",x"79"),
   940 => (x"00",x"76",x"00",x"05"),
   941 => (x"00",x"0d",x"00",x"07"),
   942 => (x"00",x"1e",x"00",x"0d"),
   943 => (x"00",x"29",x"00",x"06"),
   944 => (x"04",x"14",x"00",x"00"),
   945 => (x"00",x"15",x"00",x"00"),
   946 => (x"40",x"00",x"00",x"00"),
   947 => (x"40",x"00",x"00",x"00"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

