library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"4a1387e7",
     1 => x"87f5059a",
     2 => x"1e87dafe",
     3 => x"bfd5cdc3",
     4 => x"d5cdc349",
     5 => x"78a1c148",
     6 => x"a9b7c0c4",
     7 => x"ff87db03",
     8 => x"cdc348d4",
     9 => x"c378bfd9",
    10 => x"49bfd5cd",
    11 => x"48d5cdc3",
    12 => x"c478a1c1",
    13 => x"04a9b7c0",
    14 => x"d0ff87e5",
    15 => x"c378c848",
    16 => x"c048e1cd",
    17 => x"004f2678",
    18 => x"00000000",
    19 => x"00000000",
    20 => x"5f5f0000",
    21 => x"00000000",
    22 => x"03000303",
    23 => x"14000003",
    24 => x"7f147f7f",
    25 => x"0000147f",
    26 => x"6b6b2e24",
    27 => x"4c00123a",
    28 => x"6c18366a",
    29 => x"30003256",
    30 => x"77594f7e",
    31 => x"0040683a",
    32 => x"03070400",
    33 => x"00000000",
    34 => x"633e1c00",
    35 => x"00000041",
    36 => x"3e634100",
    37 => x"0800001c",
    38 => x"1c1c3e2a",
    39 => x"00082a3e",
    40 => x"3e3e0808",
    41 => x"00000808",
    42 => x"60e08000",
    43 => x"00000000",
    44 => x"08080808",
    45 => x"00000808",
    46 => x"60600000",
    47 => x"40000000",
    48 => x"0c183060",
    49 => x"00010306",
    50 => x"4d597f3e",
    51 => x"00003e7f",
    52 => x"7f7f0604",
    53 => x"00000000",
    54 => x"59716342",
    55 => x"0000464f",
    56 => x"49496322",
    57 => x"1800367f",
    58 => x"7f13161c",
    59 => x"0000107f",
    60 => x"45456727",
    61 => x"0000397d",
    62 => x"494b7e3c",
    63 => x"00003079",
    64 => x"79710101",
    65 => x"0000070f",
    66 => x"49497f36",
    67 => x"0000367f",
    68 => x"69494f06",
    69 => x"00001e3f",
    70 => x"66660000",
    71 => x"00000000",
    72 => x"66e68000",
    73 => x"00000000",
    74 => x"14140808",
    75 => x"00002222",
    76 => x"14141414",
    77 => x"00001414",
    78 => x"14142222",
    79 => x"00000808",
    80 => x"59510302",
    81 => x"3e00060f",
    82 => x"555d417f",
    83 => x"00001e1f",
    84 => x"09097f7e",
    85 => x"00007e7f",
    86 => x"49497f7f",
    87 => x"0000367f",
    88 => x"41633e1c",
    89 => x"00004141",
    90 => x"63417f7f",
    91 => x"00001c3e",
    92 => x"49497f7f",
    93 => x"00004141",
    94 => x"09097f7f",
    95 => x"00000101",
    96 => x"49417f3e",
    97 => x"00007a7b",
    98 => x"08087f7f",
    99 => x"00007f7f",
   100 => x"7f7f4100",
   101 => x"00000041",
   102 => x"40406020",
   103 => x"7f003f7f",
   104 => x"361c087f",
   105 => x"00004163",
   106 => x"40407f7f",
   107 => x"7f004040",
   108 => x"060c067f",
   109 => x"7f007f7f",
   110 => x"180c067f",
   111 => x"00007f7f",
   112 => x"41417f3e",
   113 => x"00003e7f",
   114 => x"09097f7f",
   115 => x"3e00060f",
   116 => x"7f61417f",
   117 => x"0000407e",
   118 => x"19097f7f",
   119 => x"0000667f",
   120 => x"594d6f26",
   121 => x"0000327b",
   122 => x"7f7f0101",
   123 => x"00000101",
   124 => x"40407f3f",
   125 => x"00003f7f",
   126 => x"70703f0f",
   127 => x"7f000f3f",
   128 => x"3018307f",
   129 => x"41007f7f",
   130 => x"1c1c3663",
   131 => x"01416336",
   132 => x"7c7c0603",
   133 => x"61010306",
   134 => x"474d5971",
   135 => x"00004143",
   136 => x"417f7f00",
   137 => x"01000041",
   138 => x"180c0603",
   139 => x"00406030",
   140 => x"7f414100",
   141 => x"0800007f",
   142 => x"0603060c",
   143 => x"8000080c",
   144 => x"80808080",
   145 => x"00008080",
   146 => x"07030000",
   147 => x"00000004",
   148 => x"54547420",
   149 => x"0000787c",
   150 => x"44447f7f",
   151 => x"0000387c",
   152 => x"44447c38",
   153 => x"00000044",
   154 => x"44447c38",
   155 => x"00007f7f",
   156 => x"54547c38",
   157 => x"0000185c",
   158 => x"057f7e04",
   159 => x"00000005",
   160 => x"a4a4bc18",
   161 => x"00007cfc",
   162 => x"04047f7f",
   163 => x"0000787c",
   164 => x"7d3d0000",
   165 => x"00000040",
   166 => x"fd808080",
   167 => x"0000007d",
   168 => x"38107f7f",
   169 => x"0000446c",
   170 => x"7f3f0000",
   171 => x"7c000040",
   172 => x"0c180c7c",
   173 => x"0000787c",
   174 => x"04047c7c",
   175 => x"0000787c",
   176 => x"44447c38",
   177 => x"0000387c",
   178 => x"2424fcfc",
   179 => x"0000183c",
   180 => x"24243c18",
   181 => x"0000fcfc",
   182 => x"04047c7c",
   183 => x"0000080c",
   184 => x"54545c48",
   185 => x"00002074",
   186 => x"447f3f04",
   187 => x"00000044",
   188 => x"40407c3c",
   189 => x"00007c7c",
   190 => x"60603c1c",
   191 => x"3c001c3c",
   192 => x"6030607c",
   193 => x"44003c7c",
   194 => x"3810386c",
   195 => x"0000446c",
   196 => x"60e0bc1c",
   197 => x"00001c3c",
   198 => x"5c746444",
   199 => x"0000444c",
   200 => x"773e0808",
   201 => x"00004141",
   202 => x"7f7f0000",
   203 => x"00000000",
   204 => x"3e774141",
   205 => x"02000808",
   206 => x"02030101",
   207 => x"7f000102",
   208 => x"7f7f7f7f",
   209 => x"08007f7f",
   210 => x"3e1c1c08",
   211 => x"7f7f7f3e",
   212 => x"1c3e3e7f",
   213 => x"0008081c",
   214 => x"7c7c1810",
   215 => x"00001018",
   216 => x"7c7c3010",
   217 => x"10001030",
   218 => x"78606030",
   219 => x"4200061e",
   220 => x"3c183c66",
   221 => x"78004266",
   222 => x"c6c26a38",
   223 => x"6000386c",
   224 => x"00600000",
   225 => x"0e006000",
   226 => x"5d5c5b5e",
   227 => x"4c711e0e",
   228 => x"bff2cdc3",
   229 => x"c04bc04d",
   230 => x"02ab741e",
   231 => x"a6c487c7",
   232 => x"c578c048",
   233 => x"48a6c487",
   234 => x"66c478c1",
   235 => x"ee49731e",
   236 => x"86c887df",
   237 => x"ef49e0c0",
   238 => x"a5c487ef",
   239 => x"f0496a4a",
   240 => x"c6f187f0",
   241 => x"c185cb87",
   242 => x"abb7c883",
   243 => x"87c7ff04",
   244 => x"264d2626",
   245 => x"264b264c",
   246 => x"4a711e4f",
   247 => x"5af6cdc3",
   248 => x"48f6cdc3",
   249 => x"fe4978c7",
   250 => x"4f2687dd",
   251 => x"711e731e",
   252 => x"aab7c04a",
   253 => x"c287d303",
   254 => x"05bfc2e0",
   255 => x"4bc187c4",
   256 => x"4bc087c2",
   257 => x"5bc6e0c2",
   258 => x"e0c287c4",
   259 => x"e0c25ac6",
   260 => x"c14abfc2",
   261 => x"a2c0c19a",
   262 => x"87e8ec49",
   263 => x"bfeadfc2",
   264 => x"c2e0c249",
   265 => x"48fcb1bf",
   266 => x"e8fe7871",
   267 => x"4a711e87",
   268 => x"721e66c4",
   269 => x"dbdfff49",
   270 => x"4f262687",
   271 => x"c2e0c21e",
   272 => x"e2c049bf",
   273 => x"cdc387f0",
   274 => x"bfe848ea",
   275 => x"e6cdc378",
   276 => x"78bfec48",
   277 => x"bfeacdc3",
   278 => x"ffc3494a",
   279 => x"2ab7c899",
   280 => x"b0714872",
   281 => x"58f2cdc3",
   282 => x"5e0e4f26",
   283 => x"0e5d5c5b",
   284 => x"c7ff4b71",
   285 => x"e5cdc387",
   286 => x"7350c048",
   287 => x"e8dbff49",
   288 => x"4c497087",
   289 => x"eecb9cc2",
   290 => x"87fecd49",
   291 => x"c34d4970",
   292 => x"bf97e5cd",
   293 => x"87e4c105",
   294 => x"c34966d0",
   295 => x"99bfeecd",
   296 => x"d487d705",
   297 => x"cdc34966",
   298 => x"0599bfe6",
   299 => x"497387cc",
   300 => x"87f5daff",
   301 => x"c1029870",
   302 => x"4cc187c2",
   303 => x"7587fdfd",
   304 => x"87d2cd49",
   305 => x"c6029870",
   306 => x"e5cdc387",
   307 => x"c350c148",
   308 => x"bf97e5cd",
   309 => x"87e4c005",
   310 => x"bfeecdc3",
   311 => x"9966d049",
   312 => x"87d6ff05",
   313 => x"bfe6cdc3",
   314 => x"9966d449",
   315 => x"87caff05",
   316 => x"d9ff4973",
   317 => x"987087f3",
   318 => x"87fefe05",
   319 => x"d0fb4874",
   320 => x"5b5e0e87",
   321 => x"f80e5d5c",
   322 => x"4c4dc086",
   323 => x"c47ebfec",
   324 => x"cdc348a6",
   325 => x"c078bff2",
   326 => x"f7c11e1e",
   327 => x"87cafd49",
   328 => x"987086c8",
   329 => x"87f3c002",
   330 => x"bfeadfc2",
   331 => x"c187c405",
   332 => x"c087c27e",
   333 => x"eadfc27e",
   334 => x"ca786e48",
   335 => x"66c41efc",
   336 => x"c487c902",
   337 => x"dec248a6",
   338 => x"87c778c1",
   339 => x"c248a6c4",
   340 => x"c478ccde",
   341 => x"ffc84966",
   342 => x"c186c487",
   343 => x"c71ec01e",
   344 => x"87c6fc49",
   345 => x"987086c8",
   346 => x"ff87ce02",
   347 => x"87fcf949",
   348 => x"ff49dac1",
   349 => x"c187f2d7",
   350 => x"e5cdc34d",
   351 => x"c302bf97",
   352 => x"87e4cf87",
   353 => x"bfeacdc3",
   354 => x"c2e0c24b",
   355 => x"e4c105bf",
   356 => x"eadfc287",
   357 => x"f1c002bf",
   358 => x"48a6c487",
   359 => x"78c0c0c8",
   360 => x"7eeedfc2",
   361 => x"49bf976e",
   362 => x"80c1486e",
   363 => x"ff717e70",
   364 => x"7087f6d6",
   365 => x"87c30298",
   366 => x"c4b366c4",
   367 => x"b7c14866",
   368 => x"58a6c828",
   369 => x"ff059870",
   370 => x"fdc387da",
   371 => x"d8d6ff49",
   372 => x"49fac387",
   373 => x"87d1d6ff",
   374 => x"ffc34973",
   375 => x"c01e7199",
   376 => x"87c9f949",
   377 => x"b7c84973",
   378 => x"c11e7129",
   379 => x"87fdf849",
   380 => x"c7c686c8",
   381 => x"eecdc387",
   382 => x"029b4bbf",
   383 => x"dfc287df",
   384 => x"c849bffe",
   385 => x"987087d0",
   386 => x"87c4c005",
   387 => x"87d34bc0",
   388 => x"c749e0c2",
   389 => x"e0c287f4",
   390 => x"c6c058c2",
   391 => x"fedfc287",
   392 => x"7378c048",
   393 => x"0599c249",
   394 => x"c387cfc0",
   395 => x"d4ff49eb",
   396 => x"497087f7",
   397 => x"c00299c2",
   398 => x"4cfb87c2",
   399 => x"99c14973",
   400 => x"87cfc005",
   401 => x"ff49f4c3",
   402 => x"7087ded4",
   403 => x"0299c249",
   404 => x"fa87c2c0",
   405 => x"c849734c",
   406 => x"cfc00599",
   407 => x"49f5c387",
   408 => x"87c5d4ff",
   409 => x"99c24970",
   410 => x"87d6c002",
   411 => x"bff6cdc3",
   412 => x"87cac002",
   413 => x"c388c148",
   414 => x"c058facd",
   415 => x"4cff87c2",
   416 => x"49734dc1",
   417 => x"c00599c4",
   418 => x"f2c387cf",
   419 => x"d8d3ff49",
   420 => x"c2497087",
   421 => x"dcc00299",
   422 => x"f6cdc387",
   423 => x"c7487ebf",
   424 => x"c003a8b7",
   425 => x"486e87cb",
   426 => x"cdc380c1",
   427 => x"c2c058fa",
   428 => x"c14cfe87",
   429 => x"49fdc34d",
   430 => x"87edd2ff",
   431 => x"99c24970",
   432 => x"87d5c002",
   433 => x"bff6cdc3",
   434 => x"87c9c002",
   435 => x"48f6cdc3",
   436 => x"c2c078c0",
   437 => x"c14cfd87",
   438 => x"49fac34d",
   439 => x"87c9d2ff",
   440 => x"99c24970",
   441 => x"87d9c002",
   442 => x"bff6cdc3",
   443 => x"a8b7c748",
   444 => x"87c9c003",
   445 => x"48f6cdc3",
   446 => x"c2c078c7",
   447 => x"c14cfc87",
   448 => x"acb7c04d",
   449 => x"87d5c003",
   450 => x"c14866c4",
   451 => x"7e7080d8",
   452 => x"c002bf6e",
   453 => x"bf6e87c7",
   454 => x"7349744b",
   455 => x"c31ec00f",
   456 => x"dac11ef0",
   457 => x"87c2f549",
   458 => x"987086c8",
   459 => x"87d9c002",
   460 => x"bff6cdc3",
   461 => x"cb496e7e",
   462 => x"4a66c491",
   463 => x"026a8271",
   464 => x"6a87c6c0",
   465 => x"73496e4b",
   466 => x"029d750f",
   467 => x"c387c8c0",
   468 => x"49bff6cd",
   469 => x"c287f0f0",
   470 => x"02bfc6e0",
   471 => x"4987ddc0",
   472 => x"7087f3c2",
   473 => x"d3c00298",
   474 => x"f6cdc387",
   475 => x"d6f049bf",
   476 => x"f149c087",
   477 => x"e0c287f6",
   478 => x"78c048c6",
   479 => x"d0f18ef8",
   480 => x"796f4a87",
   481 => x"7379656b",
   482 => x"006e6f20",
   483 => x"6b796f4a",
   484 => x"20737965",
   485 => x"0066666f",
   486 => x"5c5b5e0e",
   487 => x"711e0e5d",
   488 => x"f2cdc34c",
   489 => x"cdc149bf",
   490 => x"d1c14da1",
   491 => x"747e6981",
   492 => x"87cf029c",
   493 => x"744ba5c4",
   494 => x"f2cdc37b",
   495 => x"d8f049bf",
   496 => x"747b6e87",
   497 => x"87c4059c",
   498 => x"87c24bc0",
   499 => x"49734bc1",
   500 => x"d487d9f0",
   501 => x"87c80266",
   502 => x"87eec049",
   503 => x"87c24a70",
   504 => x"e0c24ac0",
   505 => x"ef265aca",
   506 => x"000087e7",
   507 => x"12580000",
   508 => x"1b1d1411",
   509 => x"595a231c",
   510 => x"f2f59491",
   511 => x"0000f4eb",
   512 => x"00000000",
   513 => x"00000000",
   514 => x"711e0000",
   515 => x"bfc8ff4a",
   516 => x"48a17249",
   517 => x"ff1e4f26",
   518 => x"fe89bfc8",
   519 => x"c0c0c0c0",
   520 => x"c401a9c0",
   521 => x"c24ac087",
   522 => x"724ac187",
   523 => x"0e4f2648",
   524 => x"5d5c5b5e",
   525 => x"4d711e0e",
   526 => x"754bd4ff",
   527 => x"facdc31e",
   528 => x"c2c0fe49",
   529 => x"7086c487",
   530 => x"c3026e7e",
   531 => x"cec387ff",
   532 => x"754cbfc2",
   533 => x"f0d9fe49",
   534 => x"05a8de87",
   535 => x"7587ebc0",
   536 => x"f6d0ff49",
   537 => x"02987087",
   538 => x"ccc387db",
   539 => x"c01ebffd",
   540 => x"ceff49e1",
   541 => x"86c487c9",
   542 => x"48e7e5c2",
   543 => x"cdc350c0",
   544 => x"eafe49c9",
   545 => x"c348c187",
   546 => x"d0ff87c5",
   547 => x"78c5c848",
   548 => x"c07bd6c1",
   549 => x"bf976e4a",
   550 => x"c1486e7b",
   551 => x"c17e7080",
   552 => x"b7e0c082",
   553 => x"ecff04aa",
   554 => x"48d0ff87",
   555 => x"c5c878c4",
   556 => x"7bd3c178",
   557 => x"78c47bc1",
   558 => x"c1029c74",
   559 => x"fbc287fd",
   560 => x"c0c87ef6",
   561 => x"b7c08c4d",
   562 => x"87c603ac",
   563 => x"4da4c0c8",
   564 => x"c8c34cc0",
   565 => x"49bf97e7",
   566 => x"d20299d0",
   567 => x"c31ec087",
   568 => x"fe49facd",
   569 => x"c487fcc0",
   570 => x"4a497086",
   571 => x"c287efc0",
   572 => x"c31ef6fb",
   573 => x"fe49facd",
   574 => x"c487e8c0",
   575 => x"4a497086",
   576 => x"c848d0ff",
   577 => x"d4c178c5",
   578 => x"bf976e7b",
   579 => x"c1486e7b",
   580 => x"c17e7080",
   581 => x"f0ff058d",
   582 => x"48d0ff87",
   583 => x"9a7278c4",
   584 => x"87c5c005",
   585 => x"e6c048c0",
   586 => x"c31ec187",
   587 => x"fd49facd",
   588 => x"c487cffe",
   589 => x"059c7486",
   590 => x"ff87c3fe",
   591 => x"c5c848d0",
   592 => x"7bd3c178",
   593 => x"78c47bc0",
   594 => x"c2c048c1",
   595 => x"2648c087",
   596 => x"4c264d26",
   597 => x"4f264b26",
   598 => x"c44a711e",
   599 => x"87c50566",
   600 => x"cafb4972",
   601 => x"004f2687",
   602 => x"f6e6c21e",
   603 => x"b9c149bf",
   604 => x"59fae6c2",
   605 => x"c348d4ff",
   606 => x"d0ff78ff",
   607 => x"78e1c848",
   608 => x"c148d4ff",
   609 => x"7131c478",
   610 => x"48d0ff78",
   611 => x"2678e0c0",
   612 => x"e6c21e4f",
   613 => x"cdc31eea",
   614 => x"fafd49fa",
   615 => x"86c487e9",
   616 => x"c3029870",
   617 => x"87c0ff87",
   618 => x"35314f26",
   619 => x"205a484b",
   620 => x"46432020",
   621 => x"00000047",
   622 => x"fe1e0000",
   623 => x"c487f8fd",
   624 => x"c0c24966",
   625 => x"87cd0299",
   626 => x"c31ee0c3",
   627 => x"fe49d3cc",
   628 => x"c487c7ff",
   629 => x"4966c486",
   630 => x"0299c0c4",
   631 => x"f0c387cd",
   632 => x"d3ccc31e",
   633 => x"f1fefe49",
   634 => x"c486c487",
   635 => x"ffc14966",
   636 => x"c31e7199",
   637 => x"fe49d3cc",
   638 => x"fe87dffe",
   639 => x"2687f0fc",
   640 => x"5e0e4f26",
   641 => x"0e5d5c5b",
   642 => x"c086d8ff",
   643 => x"d2cec37e",
   644 => x"81c249bf",
   645 => x"1e721e71",
   646 => x"dbfd4ac6",
   647 => x"487187e8",
   648 => x"49264a26",
   649 => x"c358a6c8",
   650 => x"49bfd2ce",
   651 => x"1e7181c4",
   652 => x"4ac61e72",
   653 => x"87cedbfd",
   654 => x"4a264871",
   655 => x"a6cc4926",
   656 => x"d3f3c258",
   657 => x"cdf749bf",
   658 => x"02987087",
   659 => x"c087f9c9",
   660 => x"f5f649e0",
   661 => x"c2497087",
   662 => x"c059d7f3",
   663 => x"c449744c",
   664 => x"81d0fe91",
   665 => x"49744a69",
   666 => x"bfd2cec3",
   667 => x"c391c481",
   668 => x"7281dece",
   669 => x"d2029a79",
   670 => x"c1497287",
   671 => x"6e9a7189",
   672 => x"7080c148",
   673 => x"059a727e",
   674 => x"c187eeff",
   675 => x"acb7c284",
   676 => x"87c9ff04",
   677 => x"fcc0486e",
   678 => x"c804a8b7",
   679 => x"4cc087ea",
   680 => x"66c44a74",
   681 => x"c392c482",
   682 => x"7482dece",
   683 => x"8166c849",
   684 => x"cec391c4",
   685 => x"4a6a81de",
   686 => x"b9724969",
   687 => x"cec34b74",
   688 => x"c483bfd2",
   689 => x"decec393",
   690 => x"72ba6b83",
   691 => x"d4987148",
   692 => x"497458a6",
   693 => x"bfd2cec3",
   694 => x"c391c481",
   695 => x"6981dece",
   696 => x"48a6d47e",
   697 => x"a6d078c0",
   698 => x"4cffc35c",
   699 => x"df4966d0",
   700 => x"e2c60229",
   701 => x"4a66cc87",
   702 => x"d492e0c0",
   703 => x"ffc08266",
   704 => x"70887248",
   705 => x"48a6d84a",
   706 => x"80c478c0",
   707 => x"496e78c0",
   708 => x"e4c029df",
   709 => x"cec359a6",
   710 => x"78c148ce",
   711 => x"31c34972",
   712 => x"b1722ab7",
   713 => x"c499ffc0",
   714 => x"cef7c291",
   715 => x"6d85714d",
   716 => x"c0c4494b",
   717 => x"d70299c0",
   718 => x"66e0c087",
   719 => x"87c7c002",
   720 => x"78c080c8",
   721 => x"c387d0c5",
   722 => x"c148d6ce",
   723 => x"87c7c578",
   724 => x"0266e0c0",
   725 => x"497387d8",
   726 => x"99c0c0c2",
   727 => x"87c3c002",
   728 => x"6d2bb7d0",
   729 => x"fffffd48",
   730 => x"c07d7098",
   731 => x"cec387fa",
   732 => x"c002bfd6",
   733 => x"487387f2",
   734 => x"c028b7d0",
   735 => x"7058a6e8",
   736 => x"e3c00298",
   737 => x"dacec387",
   738 => x"e0c049bf",
   739 => x"c00299c0",
   740 => x"497087ca",
   741 => x"99c0e0c0",
   742 => x"87ccc002",
   743 => x"c0c2486d",
   744 => x"7d70b0c0",
   745 => x"4b66e4c0",
   746 => x"c0c84973",
   747 => x"c20299c0",
   748 => x"cec387c5",
   749 => x"cc4abfda",
   750 => x"c0029ac0",
   751 => x"c0c487cf",
   752 => x"d7c0028a",
   753 => x"c0028a87",
   754 => x"dcc187f8",
   755 => x"74497387",
   756 => x"c291c299",
   757 => x"1181c2f7",
   758 => x"87dbc14b",
   759 => x"99744973",
   760 => x"f7c291c2",
   761 => x"81c181c2",
   762 => x"e0c04b11",
   763 => x"c8c00266",
   764 => x"48a6dc87",
   765 => x"fec078d2",
   766 => x"48a6d887",
   767 => x"c078d2c4",
   768 => x"497387f5",
   769 => x"91c29974",
   770 => x"81c2f7c2",
   771 => x"4b1181c1",
   772 => x"0266e0c0",
   773 => x"dc87c9c0",
   774 => x"d9c148a6",
   775 => x"87d7c078",
   776 => x"c548a6d8",
   777 => x"cec078d9",
   778 => x"74497387",
   779 => x"c291c299",
   780 => x"c181c2f7",
   781 => x"c04b1181",
   782 => x"c00266e0",
   783 => x"497387db",
   784 => x"fcc7b9ff",
   785 => x"487199c0",
   786 => x"bfdacec3",
   787 => x"decec398",
   788 => x"c49b7458",
   789 => x"d3c0b3c0",
   790 => x"c7497387",
   791 => x"7199c0fc",
   792 => x"dacec348",
   793 => x"cec3b0bf",
   794 => x"9b7458de",
   795 => x"c00266d8",
   796 => x"c31e87ca",
   797 => x"f549cece",
   798 => x"86c487c0",
   799 => x"cec31e73",
   800 => x"f5f449ce",
   801 => x"dc86c487",
   802 => x"cac00266",
   803 => x"cec31e87",
   804 => x"e5f449ce",
   805 => x"d086c487",
   806 => x"30c14866",
   807 => x"6e58a6d4",
   808 => x"7030c148",
   809 => x"4866d47e",
   810 => x"a6d880c1",
   811 => x"b7e0c058",
   812 => x"f7f804a8",
   813 => x"4c66cc87",
   814 => x"b7c284c1",
   815 => x"dff704ac",
   816 => x"d2cec387",
   817 => x"7866c448",
   818 => x"268ed8ff",
   819 => x"264c264d",
   820 => x"004f264b",
   821 => x"1e000000",
   822 => x"49724ac0",
   823 => x"cec391c4",
   824 => x"79ff81de",
   825 => x"b7c682c1",
   826 => x"87ee04aa",
   827 => x"48d2cec3",
   828 => x"784040c0",
   829 => x"731e4f26",
   830 => x"f44b711e",
   831 => x"497387c4",
   832 => x"87c7f6fe",
   833 => x"0e87c8ff",
   834 => x"0e5c5b5e",
   835 => x"ff4cd4ff",
   836 => x"c5c84bd0",
   837 => x"7cd5c17b",
   838 => x"c47c66cc",
   839 => x"7bc5c87b",
   840 => x"c17cd3c1",
   841 => x"c87bc47c",
   842 => x"d4c17bc5",
   843 => x"b74ac07c",
   844 => x"87cb06a9",
   845 => x"c17cffc3",
   846 => x"aab77182",
   847 => x"c487f504",
   848 => x"7bc5c87b",
   849 => x"c07cd3c1",
   850 => x"fd7bc47c",
   851 => x"731e87ff",
   852 => x"494b711e",
   853 => x"e2c191cb",
   854 => x"82714aee",
   855 => x"97e5cdc3",
   856 => x"87d302bf",
   857 => x"1149a2ca",
   858 => x"c187cc05",
   859 => x"49c0c81e",
   860 => x"c487d4fe",
   861 => x"7387cc86",
   862 => x"f7d4fe49",
   863 => x"fe497387",
   864 => x"fd87f1d4",
   865 => x"731e87c9",
   866 => x"c24bc01e",
   867 => x"ea49e3f6",
   868 => x"987087dd",
   869 => x"c287c405",
   870 => x"fc4beff6",
   871 => x"487387f9",
   872 => x"5387ecfc",
   873 => x"32334956",
   874 => x"52202038",
   875 => x"52004d4f",
   876 => x"6c204d4f",
   877 => x"6964616f",
   878 => x"6620676e",
   879 => x"656c6961",
   880 => x"ebf40064",
   881 => x"0605f5f2",
   882 => x"0b030c04",
   883 => x"00660a83",
   884 => x"005a00fc",
   885 => x"800000da",
   886 => x"80050894",
   887 => x"80020078",
   888 => x"80030001",
   889 => x"80040009",
   890 => x"80010000",
   891 => x"00260891",
   892 => x"001d0004",
   893 => x"001c0000",
   894 => x"00250000",
   895 => x"001a000c",
   896 => x"001b0000",
   897 => x"00240000",
   898 => x"01120000",
   899 => x"002e0000",
   900 => x"002d0003",
   901 => x"00230000",
   902 => x"00360000",
   903 => x"0021000b",
   904 => x"002b0000",
   905 => x"002c0000",
   906 => x"00220000",
   907 => x"003d0000",
   908 => x"0035006c",
   909 => x"00340000",
   910 => x"003e0000",
   911 => x"00320075",
   912 => x"00330000",
   913 => x"003c0000",
   914 => x"002a006b",
   915 => x"00460000",
   916 => x"00430001",
   917 => x"003b0073",
   918 => x"00450069",
   919 => x"003a0009",
   920 => x"00420070",
   921 => x"00440072",
   922 => x"00310074",
   923 => x"00550000",
   924 => x"004d0000",
   925 => x"004b007c",
   926 => x"007b007a",
   927 => x"00490000",
   928 => x"004c0071",
   929 => x"00540084",
   930 => x"00410077",
   931 => x"00610000",
   932 => x"005b0000",
   933 => x"0052007c",
   934 => x"00f10000",
   935 => x"02590000",
   936 => x"000e0000",
   937 => x"005d005d",
   938 => x"004a0000",
   939 => x"00160079",
   940 => x"00760005",
   941 => x"000d0007",
   942 => x"001e000d",
   943 => x"00290006",
   944 => x"04140000",
   945 => x"00150000",
   946 => x"40000000",
   947 => x"40000000",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
