library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"dcfcc287",
    12 => x"48c0c84e",
    13 => x"d5c128c2",
    14 => x"ead6e5ea",
    15 => x"c1467149",
    16 => x"87f90188",
    17 => x"49dcfcc2",
    18 => x"48f4e3c2",
    19 => x"0389d089",
    20 => x"404040c0",
    21 => x"d087f640",
    22 => x"50c00581",
    23 => x"f90589c1",
    24 => x"f4e3c287",
    25 => x"f0e3c24d",
    26 => x"02ad744c",
    27 => x"0f2487c4",
    28 => x"e9c187f7",
    29 => x"e3c287d1",
    30 => x"e3c24df4",
    31 => x"ad744cf4",
    32 => x"c487c602",
    33 => x"f50f6c8c",
    34 => x"87fd0087",
    35 => x"7186fc1e",
    36 => x"49c0ff4a",
    37 => x"c0c44869",
    38 => x"487e7098",
    39 => x"87f40298",
    40 => x"fc487972",
    41 => x"0e4f268e",
    42 => x"0e5c5b5e",
    43 => x"4cc04b71",
    44 => x"029a4a13",
    45 => x"497287cd",
    46 => x"c187d1ff",
    47 => x"9a4a1384",
    48 => x"7487f305",
    49 => x"264c2648",
    50 => x"1e4f264b",
    51 => x"1e731e72",
    52 => x"02114812",
    53 => x"c34b87ca",
    54 => x"739b98df",
    55 => x"87f00288",
    56 => x"4a264b26",
    57 => x"731e4f26",
    58 => x"c11e721e",
    59 => x"87ca048b",
    60 => x"02114812",
    61 => x"028887c4",
    62 => x"4a2687f1",
    63 => x"4f264b26",
    64 => x"8148731e",
    65 => x"c502a973",
    66 => x"05531287",
    67 => x"4f2687f6",
    68 => x"711e731e",
    69 => x"4b66c84a",
    70 => x"718bc149",
    71 => x"87cf0299",
    72 => x"d4ff4812",
    73 => x"49737808",
    74 => x"99718bc1",
    75 => x"2687f105",
    76 => x"0e4f264b",
    77 => x"0e5c5b5e",
    78 => x"d4ff4a71",
    79 => x"4b66cc4c",
    80 => x"718bc149",
    81 => x"87ce0299",
    82 => x"6c7cffc3",
    83 => x"c1497352",
    84 => x"0599718b",
    85 => x"4c2687f2",
    86 => x"4f264b26",
    87 => x"ff1e731e",
    88 => x"ffc34bd4",
    89 => x"c34a6b7b",
    90 => x"496b7bff",
    91 => x"b17232c8",
    92 => x"6b7bffc3",
    93 => x"7131c84a",
    94 => x"7bffc3b2",
    95 => x"32c8496b",
    96 => x"4871b172",
    97 => x"4f264b26",
    98 => x"5c5b5e0e",
    99 => x"4d710e5d",
   100 => x"754cd4ff",
   101 => x"98ffc348",
   102 => x"e3c27c70",
   103 => x"c805bff4",
   104 => x"4866d087",
   105 => x"a6d430c9",
   106 => x"4966d058",
   107 => x"487129d8",
   108 => x"7098ffc3",
   109 => x"4966d07c",
   110 => x"487129d0",
   111 => x"7098ffc3",
   112 => x"4966d07c",
   113 => x"487129c8",
   114 => x"7098ffc3",
   115 => x"4866d07c",
   116 => x"7098ffc3",
   117 => x"d049757c",
   118 => x"c3487129",
   119 => x"7c7098ff",
   120 => x"f0c94b6c",
   121 => x"ffc34aff",
   122 => x"87cf05ab",
   123 => x"6c7c7149",
   124 => x"028ac14b",
   125 => x"ab7187c5",
   126 => x"7387f202",
   127 => x"264d2648",
   128 => x"264b264c",
   129 => x"49c01e4f",
   130 => x"c348d4ff",
   131 => x"81c178ff",
   132 => x"a9b7c8c3",
   133 => x"2687f104",
   134 => x"5b5e0e4f",
   135 => x"c00e5d5c",
   136 => x"f7c1f0ff",
   137 => x"c0c0c14d",
   138 => x"4bc0c0c0",
   139 => x"c487d6ff",
   140 => x"c04cdff8",
   141 => x"fd49751e",
   142 => x"86c487ce",
   143 => x"c005a8c1",
   144 => x"d4ff87e5",
   145 => x"78ffc348",
   146 => x"e1c01e73",
   147 => x"49e9c1f0",
   148 => x"c487f5fc",
   149 => x"05987086",
   150 => x"d4ff87ca",
   151 => x"78ffc348",
   152 => x"87cb48c1",
   153 => x"c187defe",
   154 => x"c6ff058c",
   155 => x"2648c087",
   156 => x"264c264d",
   157 => x"0e4f264b",
   158 => x"0e5c5b5e",
   159 => x"c1f0ffc0",
   160 => x"d4ff4cc1",
   161 => x"78ffc348",
   162 => x"f849fcca",
   163 => x"4bd387d9",
   164 => x"49741ec0",
   165 => x"c487f1fb",
   166 => x"05987086",
   167 => x"d4ff87ca",
   168 => x"78ffc348",
   169 => x"87cb48c1",
   170 => x"c187dafd",
   171 => x"dfff058b",
   172 => x"2648c087",
   173 => x"264b264c",
   174 => x"0000004f",
   175 => x"00444d43",
   176 => x"43484453",
   177 => x"69616620",
   178 => x"000a216c",
   179 => x"52524549",
   180 => x"00000000",
   181 => x"00495053",
   182 => x"74697257",
   183 => x"61662065",
   184 => x"64656c69",
   185 => x"5e0e000a",
   186 => x"0e5d5c5b",
   187 => x"ff4dffc3",
   188 => x"d0fc4bd4",
   189 => x"1eeac687",
   190 => x"c1f0e1c0",
   191 => x"c7fa49c8",
   192 => x"c186c487",
   193 => x"87c802a8",
   194 => x"c087ecfd",
   195 => x"87e8c148",
   196 => x"7087c9f9",
   197 => x"ffffcf49",
   198 => x"a9eac699",
   199 => x"fd87c802",
   200 => x"48c087d5",
   201 => x"7587d1c1",
   202 => x"4cf1c07b",
   203 => x"7087eafb",
   204 => x"ecc00298",
   205 => x"c01ec087",
   206 => x"fac1f0ff",
   207 => x"87c8f949",
   208 => x"987086c4",
   209 => x"7587da05",
   210 => x"75496b7b",
   211 => x"757b757b",
   212 => x"c17b757b",
   213 => x"c40299c0",
   214 => x"db48c187",
   215 => x"d748c087",
   216 => x"05acc287",
   217 => x"c0cb87ca",
   218 => x"87fbf449",
   219 => x"87c848c0",
   220 => x"fe058cc1",
   221 => x"48c087f6",
   222 => x"4c264d26",
   223 => x"4f264b26",
   224 => x"5c5b5e0e",
   225 => x"d0ff0e5d",
   226 => x"d0e5c04d",
   227 => x"c24cc0c1",
   228 => x"c148f4e3",
   229 => x"49d4cb78",
   230 => x"c787ccf4",
   231 => x"f97dc24b",
   232 => x"7dc387e3",
   233 => x"49741ec0",
   234 => x"c487ddf7",
   235 => x"05a8c186",
   236 => x"c24b87c1",
   237 => x"87cb05ab",
   238 => x"f349cccb",
   239 => x"48c087e9",
   240 => x"c187f6c0",
   241 => x"d4ff058b",
   242 => x"87dafc87",
   243 => x"58f8e3c2",
   244 => x"cd059870",
   245 => x"c01ec187",
   246 => x"d0c1f0ff",
   247 => x"87e8f649",
   248 => x"d4ff86c4",
   249 => x"78ffc348",
   250 => x"c287eec4",
   251 => x"c258fce3",
   252 => x"48d4ff7d",
   253 => x"c178ffc3",
   254 => x"264d2648",
   255 => x"264b264c",
   256 => x"5b5e0e4f",
   257 => x"710e5d5c",
   258 => x"4cffc34d",
   259 => x"744bd4ff",
   260 => x"48d0ff7b",
   261 => x"7478c3c4",
   262 => x"c01e757b",
   263 => x"d8c1f0ff",
   264 => x"87e4f549",
   265 => x"987086c4",
   266 => x"cb87cb02",
   267 => x"f6f149d8",
   268 => x"c048c187",
   269 => x"7b7487ee",
   270 => x"c87bfec3",
   271 => x"66d41ec0",
   272 => x"87ccf349",
   273 => x"7b7486c4",
   274 => x"7b747b74",
   275 => x"4ae0dad8",
   276 => x"056b7b74",
   277 => x"8ac187c5",
   278 => x"7487f505",
   279 => x"48d0ff7b",
   280 => x"48c078c2",
   281 => x"4c264d26",
   282 => x"4f264b26",
   283 => x"5c5b5e0e",
   284 => x"86fc0e5d",
   285 => x"d4ff4b71",
   286 => x"c57ec04c",
   287 => x"4adfcdee",
   288 => x"6c7cffc3",
   289 => x"a8fec348",
   290 => x"87f8c005",
   291 => x"9b734d74",
   292 => x"d487cc02",
   293 => x"49731e66",
   294 => x"c487d8f2",
   295 => x"ff87d486",
   296 => x"d1c448d0",
   297 => x"4a66d478",
   298 => x"c17dffc3",
   299 => x"87f8058a",
   300 => x"c35aa6d8",
   301 => x"737c7cff",
   302 => x"87c5059b",
   303 => x"d048d0ff",
   304 => x"7e4ac178",
   305 => x"fe058ac1",
   306 => x"486e87f6",
   307 => x"4d268efc",
   308 => x"4b264c26",
   309 => x"731e4f26",
   310 => x"c04a711e",
   311 => x"48d4ff4b",
   312 => x"ff78ffc3",
   313 => x"c3c448d0",
   314 => x"48d4ff78",
   315 => x"7278ffc3",
   316 => x"f0ffc01e",
   317 => x"f249d1c1",
   318 => x"86c487ce",
   319 => x"d2059870",
   320 => x"1ec0c887",
   321 => x"fd4966cc",
   322 => x"86c487e2",
   323 => x"d0ff4b70",
   324 => x"7378c248",
   325 => x"264b2648",
   326 => x"5b5e0e4f",
   327 => x"c00e5d5c",
   328 => x"f0ffc01e",
   329 => x"f149c9c1",
   330 => x"1ed287de",
   331 => x"49c4e4c2",
   332 => x"c887f9fc",
   333 => x"c14cc086",
   334 => x"acb7d284",
   335 => x"c287f804",
   336 => x"bf97c4e4",
   337 => x"99c0c349",
   338 => x"05a9c0c1",
   339 => x"c287e7c0",
   340 => x"bf97cbe4",
   341 => x"c231d049",
   342 => x"bf97cce4",
   343 => x"7232c84a",
   344 => x"cde4c2b1",
   345 => x"b14abf97",
   346 => x"ffcf4c71",
   347 => x"c19cffff",
   348 => x"c134ca84",
   349 => x"e4c287e7",
   350 => x"49bf97cd",
   351 => x"99c631c1",
   352 => x"97cee4c2",
   353 => x"b7c74abf",
   354 => x"c2b1722a",
   355 => x"bf97c9e4",
   356 => x"9dcf4d4a",
   357 => x"97cae4c2",
   358 => x"9ac34abf",
   359 => x"e4c232ca",
   360 => x"4bbf97cb",
   361 => x"b27333c2",
   362 => x"97cce4c2",
   363 => x"c0c34bbf",
   364 => x"2bb7c69b",
   365 => x"81c2b273",
   366 => x"307148c1",
   367 => x"48c14970",
   368 => x"4d703075",
   369 => x"84c14c72",
   370 => x"c0c89471",
   371 => x"cc06adb7",
   372 => x"b734c187",
   373 => x"b7c0c82d",
   374 => x"f4ff01ad",
   375 => x"26487487",
   376 => x"264c264d",
   377 => x"0e4f264b",
   378 => x"5d5c5b5e",
   379 => x"c286fc0e",
   380 => x"c048ecec",
   381 => x"e4e4c278",
   382 => x"fb49c01e",
   383 => x"86c487d8",
   384 => x"c5059870",
   385 => x"c948c087",
   386 => x"4dc087d4",
   387 => x"48e8f1c2",
   388 => x"e5c278c1",
   389 => x"e1c04ada",
   390 => x"4bc849f4",
   391 => x"7087c7eb",
   392 => x"87c60598",
   393 => x"48e8f1c2",
   394 => x"e5c278c0",
   395 => x"e2c04af6",
   396 => x"4bc849c0",
   397 => x"7087efea",
   398 => x"87c60598",
   399 => x"48e8f1c2",
   400 => x"f1c278c0",
   401 => x"c002bfe8",
   402 => x"ebc287fe",
   403 => x"c24dbfea",
   404 => x"bf9fe2ec",
   405 => x"c5486e7e",
   406 => x"05a8ead6",
   407 => x"ebc287c7",
   408 => x"ce4dbfea",
   409 => x"ca486e87",
   410 => x"02a8d5e9",
   411 => x"48c087c5",
   412 => x"c287ebc7",
   413 => x"751ee4e4",
   414 => x"87daf949",
   415 => x"987086c4",
   416 => x"c087c505",
   417 => x"87d6c748",
   418 => x"4af6e5c2",
   419 => x"49cce2c0",
   420 => x"d1e94bc8",
   421 => x"05987087",
   422 => x"ecc287c8",
   423 => x"78c148ec",
   424 => x"e5c287d8",
   425 => x"e2c04ada",
   426 => x"4bc849d8",
   427 => x"7087f7e8",
   428 => x"c5c00298",
   429 => x"c648c087",
   430 => x"ecc287e4",
   431 => x"49bf97e2",
   432 => x"05a9d5c1",
   433 => x"c287cdc0",
   434 => x"bf97e3ec",
   435 => x"a9eac249",
   436 => x"87c5c002",
   437 => x"c5c648c0",
   438 => x"e4e4c287",
   439 => x"6e7ebf97",
   440 => x"a8e9c348",
   441 => x"87cec002",
   442 => x"ebc3486e",
   443 => x"c5c002a8",
   444 => x"c548c087",
   445 => x"e4c287e8",
   446 => x"49bf97ef",
   447 => x"ccc00599",
   448 => x"f0e4c287",
   449 => x"c249bf97",
   450 => x"c5c002a9",
   451 => x"c548c087",
   452 => x"e4c287cc",
   453 => x"48bf97f1",
   454 => x"58e8ecc2",
   455 => x"c1484c70",
   456 => x"ececc288",
   457 => x"f2e4c258",
   458 => x"7549bf97",
   459 => x"f3e4c281",
   460 => x"c84abf97",
   461 => x"7ea17232",
   462 => x"48c4f1c2",
   463 => x"e4c2786e",
   464 => x"48bf97f4",
   465 => x"58dcf1c2",
   466 => x"bfececc2",
   467 => x"87d3c202",
   468 => x"4af6e5c2",
   469 => x"49e8e1c0",
   470 => x"c9e64bc8",
   471 => x"02987087",
   472 => x"c087c5c0",
   473 => x"87f6c348",
   474 => x"bfe4ecc2",
   475 => x"d8f1c24c",
   476 => x"c9e5c25c",
   477 => x"c849bf97",
   478 => x"c8e5c231",
   479 => x"a14abf97",
   480 => x"cae5c249",
   481 => x"d04abf97",
   482 => x"49a17232",
   483 => x"97cbe5c2",
   484 => x"32d84abf",
   485 => x"c249a172",
   486 => x"c259e0f1",
   487 => x"91bfd8f1",
   488 => x"bfc4f1c2",
   489 => x"ccf1c281",
   490 => x"d1e5c259",
   491 => x"c84abf97",
   492 => x"d0e5c232",
   493 => x"a24bbf97",
   494 => x"d2e5c24a",
   495 => x"d04bbf97",
   496 => x"4aa27333",
   497 => x"97d3e5c2",
   498 => x"9bcf4bbf",
   499 => x"a27333d8",
   500 => x"d0f1c24a",
   501 => x"748ac25a",
   502 => x"d0f1c292",
   503 => x"78a17248",
   504 => x"c287c7c1",
   505 => x"bf97f6e4",
   506 => x"c231c849",
   507 => x"bf97f5e4",
   508 => x"c549a14a",
   509 => x"81ffc731",
   510 => x"f1c229c9",
   511 => x"e4c259d8",
   512 => x"4abf97fb",
   513 => x"e4c232c8",
   514 => x"4bbf97fa",
   515 => x"f1c24aa2",
   516 => x"f1c25ae0",
   517 => x"6e92bfd8",
   518 => x"d4f1c282",
   519 => x"ccf1c25a",
   520 => x"c278c048",
   521 => x"7248c8f1",
   522 => x"f1c278a1",
   523 => x"f1c248e0",
   524 => x"c278bfcc",
   525 => x"c248e4f1",
   526 => x"78bfd0f1",
   527 => x"bfececc2",
   528 => x"87c9c002",
   529 => x"30c44874",
   530 => x"c9c07e70",
   531 => x"d4f1c287",
   532 => x"30c448bf",
   533 => x"ecc27e70",
   534 => x"786e48f0",
   535 => x"8efc48c1",
   536 => x"4c264d26",
   537 => x"4f264b26",
   538 => x"33544146",
   539 => x"20202032",
   540 => x"00000000",
   541 => x"31544146",
   542 => x"20202036",
   543 => x"00000000",
   544 => x"33544146",
   545 => x"20202032",
   546 => x"00000000",
   547 => x"33544146",
   548 => x"20202032",
   549 => x"00000000",
   550 => x"31544146",
   551 => x"20202036",
   552 => x"5b5e0e00",
   553 => x"710e5d5c",
   554 => x"ececc24a",
   555 => x"87cb02bf",
   556 => x"2bc74b72",
   557 => x"ffc14d72",
   558 => x"7287c99d",
   559 => x"722bc84b",
   560 => x"9dffc34d",
   561 => x"bfc4f1c2",
   562 => x"ecf9c083",
   563 => x"d902abbf",
   564 => x"f0f9c087",
   565 => x"e4e4c25b",
   566 => x"ef49731e",
   567 => x"86c487f8",
   568 => x"c5059870",
   569 => x"c048c087",
   570 => x"ecc287e6",
   571 => x"d202bfec",
   572 => x"c4497587",
   573 => x"e4e4c291",
   574 => x"cf4c6981",
   575 => x"ffffffff",
   576 => x"7587cb9c",
   577 => x"c291c249",
   578 => x"9f81e4e4",
   579 => x"48744c69",
   580 => x"4c264d26",
   581 => x"4f264b26",
   582 => x"5c5b5e0e",
   583 => x"86f40e5d",
   584 => x"c459a6c8",
   585 => x"80c84866",
   586 => x"486e7e70",
   587 => x"c11e78c0",
   588 => x"87fdcc49",
   589 => x"4c7086c4",
   590 => x"fcc0029c",
   591 => x"f4ecc287",
   592 => x"4966dc4a",
   593 => x"87c3deff",
   594 => x"c0029870",
   595 => x"4a7487eb",
   596 => x"cb4966dc",
   597 => x"cddeff4b",
   598 => x"02987087",
   599 => x"1ec087db",
   600 => x"c4029c74",
   601 => x"c24dc087",
   602 => x"754dc187",
   603 => x"87c1cc49",
   604 => x"4c7086c4",
   605 => x"c4ff059c",
   606 => x"029c7487",
   607 => x"dc87f4c1",
   608 => x"486e49a4",
   609 => x"a4da7869",
   610 => x"4d66c449",
   611 => x"699f85c4",
   612 => x"ececc27d",
   613 => x"87d202bf",
   614 => x"9f49a4d4",
   615 => x"ffc04969",
   616 => x"487199ff",
   617 => x"7e7030d0",
   618 => x"7ec087c2",
   619 => x"6d48496e",
   620 => x"c47d7080",
   621 => x"78c04866",
   622 => x"cc4966c4",
   623 => x"c4796d81",
   624 => x"81d04966",
   625 => x"a6c879c0",
   626 => x"c878c048",
   627 => x"66c44c66",
   628 => x"7482d44a",
   629 => x"7291c849",
   630 => x"41c049a1",
   631 => x"84c1796d",
   632 => x"04acb7c6",
   633 => x"c487e7ff",
   634 => x"c4c14966",
   635 => x"c179c081",
   636 => x"c087c248",
   637 => x"268ef448",
   638 => x"264c264d",
   639 => x"0e4f264b",
   640 => x"5d5c5b5e",
   641 => x"d04c710e",
   642 => x"496c4d66",
   643 => x"c2b97585",
   644 => x"4abfe8ec",
   645 => x"9972baff",
   646 => x"c0029971",
   647 => x"a4c487e4",
   648 => x"f9496b4b",
   649 => x"7b7087fb",
   650 => x"bfe4ecc2",
   651 => x"71816c49",
   652 => x"c2b9757c",
   653 => x"4abfe8ec",
   654 => x"9972baff",
   655 => x"ff059971",
   656 => x"7c7587dc",
   657 => x"4c264d26",
   658 => x"4f264b26",
   659 => x"711e731e",
   660 => x"c8f1c24b",
   661 => x"a3c449bf",
   662 => x"c24a6a4a",
   663 => x"e4ecc28a",
   664 => x"a17292bf",
   665 => x"e8ecc249",
   666 => x"9a6b4abf",
   667 => x"c049a172",
   668 => x"c859f0f9",
   669 => x"e9711e66",
   670 => x"86c487dc",
   671 => x"c4059870",
   672 => x"c248c087",
   673 => x"2648c187",
   674 => x"1e4f264b",
   675 => x"4b711e73",
   676 => x"bfc8f1c2",
   677 => x"4aa3c449",
   678 => x"8ac24a6a",
   679 => x"bfe4ecc2",
   680 => x"49a17292",
   681 => x"bfe8ecc2",
   682 => x"729a6b4a",
   683 => x"f9c049a1",
   684 => x"66c859f0",
   685 => x"c8e5711e",
   686 => x"7086c487",
   687 => x"87c40598",
   688 => x"87c248c0",
   689 => x"4b2648c1",
   690 => x"5e0e4f26",
   691 => x"0e5d5c5b",
   692 => x"4b7186e4",
   693 => x"4866ecc0",
   694 => x"a6cc28c9",
   695 => x"e8ecc258",
   696 => x"b9ff49bf",
   697 => x"66c84871",
   698 => x"58a6d498",
   699 => x"986b4871",
   700 => x"c458a6d0",
   701 => x"a6c47ea3",
   702 => x"78bf6e48",
   703 => x"cc4866d0",
   704 => x"c605a866",
   705 => x"7b66c887",
   706 => x"d487c6c3",
   707 => x"ffc148a6",
   708 => x"ffffffff",
   709 => x"ff80c478",
   710 => x"d44ac078",
   711 => x"49724da3",
   712 => x"a17591c8",
   713 => x"4c66d049",
   714 => x"b7c08c69",
   715 => x"87cd04ac",
   716 => x"acb766d4",
   717 => x"dc87c603",
   718 => x"a6d85aa6",
   719 => x"c682c15c",
   720 => x"ff04aab7",
   721 => x"66d887d5",
   722 => x"a8b7c048",
   723 => x"d887d004",
   724 => x"91c84966",
   725 => x"2149a175",
   726 => x"69486e7b",
   727 => x"c087c978",
   728 => x"49a3cc7b",
   729 => x"7869486e",
   730 => x"6b4866c8",
   731 => x"58a6cc88",
   732 => x"bfe4ecc2",
   733 => x"7090c848",
   734 => x"4866c87e",
   735 => x"c901a86e",
   736 => x"4866c887",
   737 => x"c003a86e",
   738 => x"c4c187fd",
   739 => x"bf6e7ea3",
   740 => x"7591c849",
   741 => x"66cc49a1",
   742 => x"49bf6e79",
   743 => x"a17591c8",
   744 => x"6681c449",
   745 => x"48a6d079",
   746 => x"d078bf6e",
   747 => x"a8c54866",
   748 => x"c487c705",
   749 => x"78c048a6",
   750 => x"66d087c8",
   751 => x"c880c148",
   752 => x"486e58a6",
   753 => x"c87866c4",
   754 => x"49731e66",
   755 => x"c487f0f8",
   756 => x"e4e4c286",
   757 => x"f949731e",
   758 => x"a3d087f2",
   759 => x"66f0c049",
   760 => x"268ee079",
   761 => x"264c264d",
   762 => x"0e4f264b",
   763 => x"0e5c5b5e",
   764 => x"4bc04a71",
   765 => x"c0029a72",
   766 => x"a2da87e0",
   767 => x"4b699f49",
   768 => x"bfececc2",
   769 => x"d487cf02",
   770 => x"699f49a2",
   771 => x"ffc04c49",
   772 => x"34d09cff",
   773 => x"4cc087c2",
   774 => x"9b73b374",
   775 => x"4a87df02",
   776 => x"ecc28ac2",
   777 => x"9249bfe4",
   778 => x"bfc8f1c2",
   779 => x"c2807248",
   780 => x"7158e8f1",
   781 => x"c230c448",
   782 => x"c058f4ec",
   783 => x"f1c287e9",
   784 => x"c24bbfcc",
   785 => x"c248e4f1",
   786 => x"78bfd0f1",
   787 => x"bfececc2",
   788 => x"c287c902",
   789 => x"49bfe4ec",
   790 => x"87c731c4",
   791 => x"bfd4f1c2",
   792 => x"c231c449",
   793 => x"c259f4ec",
   794 => x"265be4f1",
   795 => x"264b264c",
   796 => x"5b5e0e4f",
   797 => x"f00e5d5c",
   798 => x"59a6c886",
   799 => x"ffffffcf",
   800 => x"7ec04cf8",
   801 => x"d80266c4",
   802 => x"e0e4c287",
   803 => x"c278c048",
   804 => x"c248d8e4",
   805 => x"78bfe4f1",
   806 => x"48dce4c2",
   807 => x"bfe0f1c2",
   808 => x"c1edc278",
   809 => x"c250c048",
   810 => x"49bff0ec",
   811 => x"bfe0e4c2",
   812 => x"03aa714a",
   813 => x"7287ccc4",
   814 => x"0599cf49",
   815 => x"c087eac0",
   816 => x"c248ecf9",
   817 => x"78bfd8e4",
   818 => x"1ee4e4c2",
   819 => x"bfd8e4c2",
   820 => x"d8e4c249",
   821 => x"78a1c148",
   822 => x"f9dfff71",
   823 => x"c086c487",
   824 => x"c248e8f9",
   825 => x"cc78e4e4",
   826 => x"e8f9c087",
   827 => x"e0c048bf",
   828 => x"ecf9c080",
   829 => x"e0e4c258",
   830 => x"80c148bf",
   831 => x"58e4e4c2",
   832 => x"000e6827",
   833 => x"bf97bf00",
   834 => x"c2029d4d",
   835 => x"e5c387e5",
   836 => x"dec202ad",
   837 => x"e8f9c087",
   838 => x"a3cb4bbf",
   839 => x"cf4c1149",
   840 => x"d2c105ac",
   841 => x"df497587",
   842 => x"cd89c199",
   843 => x"f4ecc291",
   844 => x"4aa3c181",
   845 => x"a3c35112",
   846 => x"c551124a",
   847 => x"51124aa3",
   848 => x"124aa3c7",
   849 => x"4aa3c951",
   850 => x"a3ce5112",
   851 => x"d051124a",
   852 => x"51124aa3",
   853 => x"124aa3d2",
   854 => x"4aa3d451",
   855 => x"a3d65112",
   856 => x"d851124a",
   857 => x"51124aa3",
   858 => x"124aa3dc",
   859 => x"4aa3de51",
   860 => x"7ec15112",
   861 => x"7487fcc0",
   862 => x"0599c849",
   863 => x"7487edc0",
   864 => x"0599d049",
   865 => x"e0c087d3",
   866 => x"ccc00266",
   867 => x"c0497387",
   868 => x"700f66e0",
   869 => x"d3c00298",
   870 => x"c0056e87",
   871 => x"ecc287c6",
   872 => x"50c048f4",
   873 => x"bfe8f9c0",
   874 => x"87e9c248",
   875 => x"48c1edc2",
   876 => x"c27e50c0",
   877 => x"49bff0ec",
   878 => x"bfe0e4c2",
   879 => x"04aa714a",
   880 => x"cf87f4fb",
   881 => x"f8ffffff",
   882 => x"e4f1c24c",
   883 => x"c8c005bf",
   884 => x"ececc287",
   885 => x"fac102bf",
   886 => x"dce4c287",
   887 => x"c0eb49bf",
   888 => x"e0e4c287",
   889 => x"48a6c458",
   890 => x"bfdce4c2",
   891 => x"ececc278",
   892 => x"dbc002bf",
   893 => x"4966c487",
   894 => x"a9749974",
   895 => x"87c8c002",
   896 => x"c048a6c8",
   897 => x"87e7c078",
   898 => x"c148a6c8",
   899 => x"87dfc078",
   900 => x"cf4966c4",
   901 => x"a999f8ff",
   902 => x"87c8c002",
   903 => x"c048a6cc",
   904 => x"87c5c078",
   905 => x"c148a6cc",
   906 => x"48a6c878",
   907 => x"c87866cc",
   908 => x"dec00566",
   909 => x"4966c487",
   910 => x"ecc289c2",
   911 => x"c291bfe4",
   912 => x"48bfc8f1",
   913 => x"e4c28071",
   914 => x"e4c258dc",
   915 => x"78c048e0",
   916 => x"c087d4f9",
   917 => x"ffffcf48",
   918 => x"f04cf8ff",
   919 => x"264d268e",
   920 => x"264b264c",
   921 => x"0000004f",
   922 => x"00000000",
   923 => x"ffffffff",
   924 => x"48d4ff1e",
   925 => x"6878ffc3",
   926 => x"1e4f2648",
   927 => x"c348d4ff",
   928 => x"d0ff78ff",
   929 => x"78e1c048",
   930 => x"d448d4ff",
   931 => x"1e4f2678",
   932 => x"c048d0ff",
   933 => x"4f2678e0",
   934 => x"87d4ff1e",
   935 => x"02994970",
   936 => x"fbc087c6",
   937 => x"87f105a9",
   938 => x"4f264871",
   939 => x"5c5b5e0e",
   940 => x"c04b710e",
   941 => x"87f8fe4c",
   942 => x"02994970",
   943 => x"c087f9c0",
   944 => x"c002a9ec",
   945 => x"fbc087f2",
   946 => x"ebc002a9",
   947 => x"b766cc87",
   948 => x"87c703ac",
   949 => x"c20266d0",
   950 => x"71537187",
   951 => x"87c20299",
   952 => x"cbfe84c1",
   953 => x"99497087",
   954 => x"c087cd02",
   955 => x"c702a9ec",
   956 => x"a9fbc087",
   957 => x"87d5ff05",
   958 => x"c30266d0",
   959 => x"7b97c087",
   960 => x"05a9fbc0",
   961 => x"4a7487c7",
   962 => x"c28a0ac0",
   963 => x"724a7487",
   964 => x"264c2648",
   965 => x"1e4f264b",
   966 => x"7087d5fd",
   967 => x"a9f0c049",
   968 => x"c087c904",
   969 => x"c301a9f9",
   970 => x"89f0c087",
   971 => x"04a9c1c1",
   972 => x"dac187c9",
   973 => x"87c301a9",
   974 => x"7189f7c0",
   975 => x"0e4f2648",
   976 => x"5d5c5b5e",
   977 => x"7186f80e",
   978 => x"fc7ec04c",
   979 => x"4bc087ed",
   980 => x"97e0ffc0",
   981 => x"a9c049bf",
   982 => x"fc87cf04",
   983 => x"83c187fa",
   984 => x"97e0ffc0",
   985 => x"06ab49bf",
   986 => x"ffc087f1",
   987 => x"02bf97e0",
   988 => x"fbfb87cf",
   989 => x"99497087",
   990 => x"c087c602",
   991 => x"f105a9ec",
   992 => x"fb4bc087",
   993 => x"4d7087ea",
   994 => x"c887e5fb",
   995 => x"dffb58a6",
   996 => x"c14a7087",
   997 => x"49a4c883",
   998 => x"ad496997",
   999 => x"c987da05",
  1000 => x"699749a4",
  1001 => x"a966c449",
  1002 => x"ca87ce05",
  1003 => x"699749a4",
  1004 => x"c405aa49",
  1005 => x"d07ec187",
  1006 => x"adecc087",
  1007 => x"c087c602",
  1008 => x"c405adfb",
  1009 => x"c14bc087",
  1010 => x"fe026e7e",
  1011 => x"fefa87f5",
  1012 => x"f8487387",
  1013 => x"264d268e",
  1014 => x"264b264c",
  1015 => x"0000004f",
  1016 => x"1e731e00",
  1017 => x"c84bd4ff",
  1018 => x"d0ff4a66",
  1019 => x"78c5c848",
  1020 => x"c148d4ff",
  1021 => x"7b1178d4",
  1022 => x"f9058ac1",
  1023 => x"48d0ff87",
  1024 => x"4b2678c4",
  1025 => x"5e0e4f26",
  1026 => x"0e5d5c5b",
  1027 => x"7e7186f8",
  1028 => x"f1c21e6e",
  1029 => x"ffe349f8",
  1030 => x"7086c487",
  1031 => x"e4c40298",
  1032 => x"c8edc187",
  1033 => x"496e4cbf",
  1034 => x"c887d4fc",
  1035 => x"987058a6",
  1036 => x"c487c505",
  1037 => x"78c148a6",
  1038 => x"c548d0ff",
  1039 => x"48d4ff78",
  1040 => x"c478d5c1",
  1041 => x"89c14966",
  1042 => x"edc131c6",
  1043 => x"4abf97c0",
  1044 => x"ffb07148",
  1045 => x"ff7808d4",
  1046 => x"78c448d0",
  1047 => x"97f4f1c2",
  1048 => x"99d049bf",
  1049 => x"c587dd02",
  1050 => x"48d4ff78",
  1051 => x"c078d6c1",
  1052 => x"48d4ff4a",
  1053 => x"c178ffc3",
  1054 => x"aae0c082",
  1055 => x"ff87f204",
  1056 => x"78c448d0",
  1057 => x"c348d4ff",
  1058 => x"d0ff78ff",
  1059 => x"ff78c548",
  1060 => x"d3c148d4",
  1061 => x"ff78c178",
  1062 => x"78c448d0",
  1063 => x"06acb7c0",
  1064 => x"c287cbc2",
  1065 => x"4bbfc0f2",
  1066 => x"737e748c",
  1067 => x"ddc1029b",
  1068 => x"4dc0c887",
  1069 => x"abb7c08b",
  1070 => x"c887c603",
  1071 => x"c04da3c0",
  1072 => x"f4f1c24b",
  1073 => x"d049bf97",
  1074 => x"87cf0299",
  1075 => x"f1c21ec0",
  1076 => x"f7e549f8",
  1077 => x"7086c487",
  1078 => x"c287d84c",
  1079 => x"c21ee4e4",
  1080 => x"e549f8f1",
  1081 => x"4c7087e6",
  1082 => x"e4c21e75",
  1083 => x"f0fb49e4",
  1084 => x"7486c887",
  1085 => x"87c5059c",
  1086 => x"cac148c0",
  1087 => x"c21ec187",
  1088 => x"e349f8f1",
  1089 => x"86c487f9",
  1090 => x"fe059b73",
  1091 => x"4c6e87e3",
  1092 => x"06acb7c0",
  1093 => x"f1c287d1",
  1094 => x"78c048f8",
  1095 => x"78c080d0",
  1096 => x"f2c280f4",
  1097 => x"c078bfc4",
  1098 => x"fd01acb7",
  1099 => x"d0ff87f5",
  1100 => x"ff78c548",
  1101 => x"d3c148d4",
  1102 => x"ff78c078",
  1103 => x"78c448d0",
  1104 => x"c2c048c1",
  1105 => x"f848c087",
  1106 => x"264d268e",
  1107 => x"264b264c",
  1108 => x"5b5e0e4f",
  1109 => x"fc0e5d5c",
  1110 => x"c04d7186",
  1111 => x"04ad4c4b",
  1112 => x"c087e8c0",
  1113 => x"741efffc",
  1114 => x"87c4029c",
  1115 => x"87c24ac0",
  1116 => x"49724ac1",
  1117 => x"c487faeb",
  1118 => x"c17e7086",
  1119 => x"c2056e83",
  1120 => x"c14b7587",
  1121 => x"06ab7584",
  1122 => x"6e87d8ff",
  1123 => x"268efc48",
  1124 => x"264c264d",
  1125 => x"0e4f264b",
  1126 => x"0e5c5b5e",
  1127 => x"66cc4b71",
  1128 => x"4c87d802",
  1129 => x"028cf0c0",
  1130 => x"4a7487d8",
  1131 => x"d1028ac1",
  1132 => x"cd028a87",
  1133 => x"c9028a87",
  1134 => x"7387d987",
  1135 => x"87c6f949",
  1136 => x"1e7487d2",
  1137 => x"d9c149c0",
  1138 => x"1e7487de",
  1139 => x"d9c14973",
  1140 => x"86c887d6",
  1141 => x"4b264c26",
  1142 => x"5e0e4f26",
  1143 => x"0e5d5c5b",
  1144 => x"4c7186fc",
  1145 => x"c291de49",
  1146 => x"714dd8f3",
  1147 => x"026d9785",
  1148 => x"c287dcc1",
  1149 => x"49bfc8f3",
  1150 => x"fd718174",
  1151 => x"7e7087d3",
  1152 => x"c0029848",
  1153 => x"f3c287f2",
  1154 => x"4a704bcc",
  1155 => x"fbfe49cb",
  1156 => x"4b7487ee",
  1157 => x"edc193cc",
  1158 => x"83c483cc",
  1159 => x"7bdcc9c1",
  1160 => x"c2c14974",
  1161 => x"7b7587fa",
  1162 => x"97c4edc1",
  1163 => x"c21e49bf",
  1164 => x"fd49ccf3",
  1165 => x"86c487e1",
  1166 => x"c2c14974",
  1167 => x"49c087e2",
  1168 => x"87fdc3c1",
  1169 => x"48f0f1c2",
  1170 => x"c04950c0",
  1171 => x"fc87c3e1",
  1172 => x"264d268e",
  1173 => x"264b264c",
  1174 => x"0000004f",
  1175 => x"64616f4c",
  1176 => x"2e676e69",
  1177 => x"00002e2e",
  1178 => x"61422080",
  1179 => x"00006b63",
  1180 => x"64616f4c",
  1181 => x"202e2a20",
  1182 => x"00000000",
  1183 => x"0000203a",
  1184 => x"61422080",
  1185 => x"00006b63",
  1186 => x"78452080",
  1187 => x"00007469",
  1188 => x"49204453",
  1189 => x"2e74696e",
  1190 => x"0000002e",
  1191 => x"00004b4f",
  1192 => x"544f4f42",
  1193 => x"20202020",
  1194 => x"004d4f52",
  1195 => x"711e731e",
  1196 => x"f3c2494b",
  1197 => x"7181bfc8",
  1198 => x"7087d6fa",
  1199 => x"c4029a4a",
  1200 => x"e6e44987",
  1201 => x"c8f3c287",
  1202 => x"7378c048",
  1203 => x"87fac149",
  1204 => x"4f264b26",
  1205 => x"711e731e",
  1206 => x"4aa3c44b",
  1207 => x"87d0c102",
  1208 => x"dc028ac1",
  1209 => x"c0028a87",
  1210 => x"058a87f2",
  1211 => x"c287d3c1",
  1212 => x"02bfc8f3",
  1213 => x"4887cbc1",
  1214 => x"f3c288c1",
  1215 => x"c1c158cc",
  1216 => x"c8f3c287",
  1217 => x"89c649bf",
  1218 => x"59ccf3c2",
  1219 => x"03a9b7c0",
  1220 => x"c287efc0",
  1221 => x"c048c8f3",
  1222 => x"87e6c078",
  1223 => x"bfc4f3c2",
  1224 => x"c287df02",
  1225 => x"48bfc8f3",
  1226 => x"f3c280c1",
  1227 => x"87d258cc",
  1228 => x"bfc4f3c2",
  1229 => x"c287cb02",
  1230 => x"48bfc8f3",
  1231 => x"f3c280c6",
  1232 => x"497358cc",
  1233 => x"4b2687c4",
  1234 => x"5e0e4f26",
  1235 => x"0e5d5c5b",
  1236 => x"a6d086f0",
  1237 => x"e4e4c259",
  1238 => x"c24cc04d",
  1239 => x"c148c4f3",
  1240 => x"48a6c878",
  1241 => x"7e7578c0",
  1242 => x"bfc8f3c2",
  1243 => x"06a8c048",
  1244 => x"c887c0c1",
  1245 => x"7e755ca6",
  1246 => x"48e4e4c2",
  1247 => x"f2c00298",
  1248 => x"4d66c487",
  1249 => x"1efffcc0",
  1250 => x"c40266cc",
  1251 => x"c24cc087",
  1252 => x"744cc187",
  1253 => x"87d9e349",
  1254 => x"7e7086c4",
  1255 => x"66c885c1",
  1256 => x"cc80c148",
  1257 => x"f3c258a6",
  1258 => x"03adbfc8",
  1259 => x"056e87c5",
  1260 => x"6e87d1ff",
  1261 => x"754cc04d",
  1262 => x"dcc3029d",
  1263 => x"fffcc087",
  1264 => x"0266cc1e",
  1265 => x"a6c887c7",
  1266 => x"c578c048",
  1267 => x"48a6c887",
  1268 => x"66c878c1",
  1269 => x"87d9e249",
  1270 => x"7e7086c4",
  1271 => x"c2029848",
  1272 => x"cb4987e4",
  1273 => x"49699781",
  1274 => x"c10299d0",
  1275 => x"497487d4",
  1276 => x"edc191cc",
  1277 => x"cac181cc",
  1278 => x"81c879ec",
  1279 => x"7451ffc3",
  1280 => x"c291de49",
  1281 => x"714dd8f3",
  1282 => x"97c1c285",
  1283 => x"49a5c17d",
  1284 => x"c251e0c0",
  1285 => x"bf97f4ec",
  1286 => x"c187d202",
  1287 => x"4ba5c284",
  1288 => x"4af4ecc2",
  1289 => x"f3fe49db",
  1290 => x"d9c187d6",
  1291 => x"49a5cd87",
  1292 => x"84c151c0",
  1293 => x"6e4ba5c2",
  1294 => x"fe49cb4a",
  1295 => x"c187c1f3",
  1296 => x"497487c4",
  1297 => x"edc191cc",
  1298 => x"c7c181cc",
  1299 => x"ecc279da",
  1300 => x"02bf97f4",
  1301 => x"497487d8",
  1302 => x"84c191de",
  1303 => x"4bd8f3c2",
  1304 => x"ecc28371",
  1305 => x"49dd4af4",
  1306 => x"87d4f2fe",
  1307 => x"4b7487d8",
  1308 => x"f3c293de",
  1309 => x"a3cb83d8",
  1310 => x"c151c049",
  1311 => x"4a6e7384",
  1312 => x"f1fe49cb",
  1313 => x"66c887fa",
  1314 => x"cc80c148",
  1315 => x"acc758a6",
  1316 => x"87c5c003",
  1317 => x"e4fc056e",
  1318 => x"03acc787",
  1319 => x"c287e4c0",
  1320 => x"c048c4f3",
  1321 => x"cc497478",
  1322 => x"ccedc191",
  1323 => x"dac7c181",
  1324 => x"de497479",
  1325 => x"d8f3c291",
  1326 => x"c151c081",
  1327 => x"04acc784",
  1328 => x"c187dcff",
  1329 => x"c048e8ee",
  1330 => x"c180f750",
  1331 => x"c140f0d4",
  1332 => x"c878e8c9",
  1333 => x"d4cbc180",
  1334 => x"4966cc78",
  1335 => x"87c0f8c0",
  1336 => x"4d268ef0",
  1337 => x"4b264c26",
  1338 => x"731e4f26",
  1339 => x"494b711e",
  1340 => x"edc191cc",
  1341 => x"a1c881cc",
  1342 => x"c0edc14a",
  1343 => x"c9501248",
  1344 => x"ffc04aa1",
  1345 => x"501248e0",
  1346 => x"edc181ca",
  1347 => x"501148c4",
  1348 => x"97c4edc1",
  1349 => x"c01e49bf",
  1350 => x"87fbf149",
  1351 => x"e9f84973",
  1352 => x"268efc87",
  1353 => x"1e4f264b",
  1354 => x"f8c049c0",
  1355 => x"4f2687d3",
  1356 => x"494a711e",
  1357 => x"edc191cc",
  1358 => x"81c881cc",
  1359 => x"48f0f1c2",
  1360 => x"f0c05011",
  1361 => x"edfe49a2",
  1362 => x"49c087c2",
  1363 => x"2687c3d5",
  1364 => x"d4ff1e4f",
  1365 => x"7affc34a",
  1366 => x"c048d0ff",
  1367 => x"7ade78e1",
  1368 => x"c8487a71",
  1369 => x"7a7028b7",
  1370 => x"b7d04871",
  1371 => x"717a7028",
  1372 => x"28b7d848",
  1373 => x"d0ff7a70",
  1374 => x"78e0c048",
  1375 => x"5e0e4f26",
  1376 => x"0e5d5c5b",
  1377 => x"4d7186f4",
  1378 => x"c191cc49",
  1379 => x"c881cced",
  1380 => x"a1ca4aa1",
  1381 => x"48a6c47e",
  1382 => x"bfecf1c2",
  1383 => x"bf976e78",
  1384 => x"4c66c44b",
  1385 => x"48122c73",
  1386 => x"7058a6cc",
  1387 => x"c984c19c",
  1388 => x"49699781",
  1389 => x"c204acb7",
  1390 => x"6e4cc087",
  1391 => x"c84abf97",
  1392 => x"31724966",
  1393 => x"66c4b9ff",
  1394 => x"72487499",
  1395 => x"b14a7030",
  1396 => x"59f0f1c2",
  1397 => x"87f9fd71",
  1398 => x"f3c21ec7",
  1399 => x"c11ebfc0",
  1400 => x"c21ecced",
  1401 => x"bf97f0f1",
  1402 => x"87f4c149",
  1403 => x"f3c04975",
  1404 => x"8ee887ee",
  1405 => x"4c264d26",
  1406 => x"4f264b26",
  1407 => x"711e731e",
  1408 => x"f9fd494b",
  1409 => x"fd497387",
  1410 => x"4b2687f4",
  1411 => x"731e4f26",
  1412 => x"c24b711e",
  1413 => x"d6024aa3",
  1414 => x"058ac187",
  1415 => x"c287e2c0",
  1416 => x"02bfc0f3",
  1417 => x"c14887db",
  1418 => x"c4f3c288",
  1419 => x"c287d258",
  1420 => x"02bfc4f3",
  1421 => x"f3c287cb",
  1422 => x"c148bfc0",
  1423 => x"c4f3c280",
  1424 => x"c21ec758",
  1425 => x"1ebfc0f3",
  1426 => x"1eccedc1",
  1427 => x"97f0f1c2",
  1428 => x"87cc49bf",
  1429 => x"f2c04973",
  1430 => x"8ef487c6",
  1431 => x"4f264b26",
  1432 => x"5c5b5e0e",
  1433 => x"ccff0e5d",
  1434 => x"a6e8c086",
  1435 => x"48a6cc59",
  1436 => x"80c478c0",
  1437 => x"80c478c0",
  1438 => x"80c478c0",
  1439 => x"7866c8c1",
  1440 => x"78c180c4",
  1441 => x"78c180c4",
  1442 => x"48c4f3c2",
  1443 => x"dfff78c1",
  1444 => x"c3e087e9",
  1445 => x"d7dfff87",
  1446 => x"c04d7087",
  1447 => x"c102adfb",
  1448 => x"e4c087f3",
  1449 => x"e8c10566",
  1450 => x"66c4c187",
  1451 => x"6a82c44a",
  1452 => x"f0c9c17e",
  1453 => x"20496e48",
  1454 => x"10412041",
  1455 => x"66c4c151",
  1456 => x"ead3c148",
  1457 => x"c7496a78",
  1458 => x"c1517581",
  1459 => x"c84966c4",
  1460 => x"dc51c181",
  1461 => x"78c248a6",
  1462 => x"4966c4c1",
  1463 => x"51c081c9",
  1464 => x"4966c4c1",
  1465 => x"51c081ca",
  1466 => x"1ed81ec1",
  1467 => x"81c8496a",
  1468 => x"87f8deff",
  1469 => x"c8c186c8",
  1470 => x"a8c04866",
  1471 => x"d487c701",
  1472 => x"78c148a6",
  1473 => x"c8c187cf",
  1474 => x"88c14866",
  1475 => x"c458a6dc",
  1476 => x"c3deff87",
  1477 => x"029d7587",
  1478 => x"d487f1cb",
  1479 => x"ccc14866",
  1480 => x"cb03a866",
  1481 => x"7ec087e6",
  1482 => x"87c4ddff",
  1483 => x"c1484d70",
  1484 => x"a6c888c6",
  1485 => x"02987058",
  1486 => x"4887d6c1",
  1487 => x"a6c888c9",
  1488 => x"02987058",
  1489 => x"4887d7c5",
  1490 => x"a6c888c1",
  1491 => x"02987058",
  1492 => x"4887f8c2",
  1493 => x"a6c888c3",
  1494 => x"02987058",
  1495 => x"c14887cf",
  1496 => x"58a6c888",
  1497 => x"c4029870",
  1498 => x"fec987f4",
  1499 => x"7ef0c087",
  1500 => x"87fcdbff",
  1501 => x"ecc04d70",
  1502 => x"87c202ad",
  1503 => x"ecc07e75",
  1504 => x"87cd02ad",
  1505 => x"87e8dbff",
  1506 => x"ecc04d70",
  1507 => x"f3ff05ad",
  1508 => x"66e4c087",
  1509 => x"87eac105",
  1510 => x"02adecc0",
  1511 => x"dbff87c4",
  1512 => x"1ec087ce",
  1513 => x"66dc1eca",
  1514 => x"c193cc4b",
  1515 => x"c48366cc",
  1516 => x"496c4ca3",
  1517 => x"87f4dbff",
  1518 => x"1ede1ec1",
  1519 => x"dbff496c",
  1520 => x"86d087ea",
  1521 => x"7bead3c1",
  1522 => x"dc49a3c8",
  1523 => x"a3c95166",
  1524 => x"66e0c049",
  1525 => x"49a3ca51",
  1526 => x"66dc516e",
  1527 => x"c080c148",
  1528 => x"d458a6e0",
  1529 => x"66d84866",
  1530 => x"87cb04a8",
  1531 => x"c14866d4",
  1532 => x"58a6d880",
  1533 => x"d887fac7",
  1534 => x"88c14866",
  1535 => x"c758a6dc",
  1536 => x"daff87ef",
  1537 => x"4d7087d2",
  1538 => x"ff87e6c7",
  1539 => x"d087c8dc",
  1540 => x"66d058a6",
  1541 => x"87c606a8",
  1542 => x"cc48a6d0",
  1543 => x"dbff7866",
  1544 => x"ecc087f5",
  1545 => x"f5c105a8",
  1546 => x"66e4c087",
  1547 => x"87e5c105",
  1548 => x"cc4966d4",
  1549 => x"66c4c191",
  1550 => x"4aa1c481",
  1551 => x"a1c84c6a",
  1552 => x"5266cc4a",
  1553 => x"79f0d4c1",
  1554 => x"87e4d8ff",
  1555 => x"029d4d70",
  1556 => x"fbc087da",
  1557 => x"87d402ad",
  1558 => x"d8ff5475",
  1559 => x"4d7087d2",
  1560 => x"c7c0029d",
  1561 => x"adfbc087",
  1562 => x"87ecff05",
  1563 => x"c254e0c0",
  1564 => x"97c054c1",
  1565 => x"4866d47c",
  1566 => x"04a866d8",
  1567 => x"d487cbc0",
  1568 => x"80c14866",
  1569 => x"c558a6d8",
  1570 => x"66d887e7",
  1571 => x"dc88c148",
  1572 => x"dcc558a6",
  1573 => x"ffd7ff87",
  1574 => x"c54d7087",
  1575 => x"66cc87d3",
  1576 => x"66e4c048",
  1577 => x"f4c405a8",
  1578 => x"a6e8c087",
  1579 => x"ff78c048",
  1580 => x"7087e4d9",
  1581 => x"ded9ff7e",
  1582 => x"a6f0c087",
  1583 => x"a8ecc058",
  1584 => x"87c7c005",
  1585 => x"786e48a6",
  1586 => x"ff87c4c0",
  1587 => x"d487e1d6",
  1588 => x"91cc4966",
  1589 => x"4866c4c1",
  1590 => x"a6c88071",
  1591 => x"4a66c458",
  1592 => x"66c482c8",
  1593 => x"6e81ca49",
  1594 => x"66ecc051",
  1595 => x"6e81c149",
  1596 => x"7148c189",
  1597 => x"c1497030",
  1598 => x"7a977189",
  1599 => x"bfecf1c2",
  1600 => x"97296e49",
  1601 => x"71484a6a",
  1602 => x"a6f4c098",
  1603 => x"4866c458",
  1604 => x"a6cc80c4",
  1605 => x"bf66c858",
  1606 => x"66e4c04c",
  1607 => x"a866cc48",
  1608 => x"87c5c002",
  1609 => x"c2c07ec0",
  1610 => x"6e7ec187",
  1611 => x"1ee0c01e",
  1612 => x"d5ff4974",
  1613 => x"86c887f6",
  1614 => x"b7c04d70",
  1615 => x"d4c106ad",
  1616 => x"c8847587",
  1617 => x"c049bf66",
  1618 => x"897481e0",
  1619 => x"fcc9c14b",
  1620 => x"defe714a",
  1621 => x"84c287ea",
  1622 => x"e8c07e74",
  1623 => x"80c14866",
  1624 => x"58a6ecc0",
  1625 => x"4966f0c0",
  1626 => x"a97081c1",
  1627 => x"87c5c002",
  1628 => x"c2c04cc0",
  1629 => x"744cc187",
  1630 => x"bf66cc1e",
  1631 => x"81e0c049",
  1632 => x"718966c4",
  1633 => x"4966c81e",
  1634 => x"87e0d4ff",
  1635 => x"b7c086c8",
  1636 => x"c5ff01a8",
  1637 => x"66e8c087",
  1638 => x"87d3c002",
  1639 => x"c94966c4",
  1640 => x"66e8c081",
  1641 => x"4866c451",
  1642 => x"78fed5c1",
  1643 => x"c487cec0",
  1644 => x"81c94966",
  1645 => x"66c451c2",
  1646 => x"fcd7c148",
  1647 => x"4866d478",
  1648 => x"04a866d8",
  1649 => x"d487cbc0",
  1650 => x"80c14866",
  1651 => x"c058a6d8",
  1652 => x"66d887d1",
  1653 => x"dc88c148",
  1654 => x"c6c058a6",
  1655 => x"f7d2ff87",
  1656 => x"cc4d7087",
  1657 => x"78c048a6",
  1658 => x"ff87c6c0",
  1659 => x"7087e9d2",
  1660 => x"66e0c04d",
  1661 => x"c080c148",
  1662 => x"7558a6e4",
  1663 => x"cbc0029d",
  1664 => x"4866d487",
  1665 => x"a866ccc1",
  1666 => x"87daf404",
  1667 => x"c74866d4",
  1668 => x"e1c003a8",
  1669 => x"4c66d487",
  1670 => x"48c4f3c2",
  1671 => x"497478c0",
  1672 => x"c4c191cc",
  1673 => x"a1c48166",
  1674 => x"c04a6a4a",
  1675 => x"84c17952",
  1676 => x"ff04acc7",
  1677 => x"e4c087e2",
  1678 => x"e2c00266",
  1679 => x"66c4c187",
  1680 => x"81d4c149",
  1681 => x"4a66c4c1",
  1682 => x"c082dcc1",
  1683 => x"f0d4c152",
  1684 => x"66c4c179",
  1685 => x"81d8c149",
  1686 => x"79c0cac1",
  1687 => x"c187d6c0",
  1688 => x"c14966c4",
  1689 => x"c4c181d4",
  1690 => x"d8c14a66",
  1691 => x"c8cac182",
  1692 => x"e7d4c17a",
  1693 => x"66c4c179",
  1694 => x"81e0c149",
  1695 => x"79ced8c1",
  1696 => x"87cbd0ff",
  1697 => x"ff4866d0",
  1698 => x"4d268ecc",
  1699 => x"4b264c26",
  1700 => x"c71e4f26",
  1701 => x"c0f3c21e",
  1702 => x"edc11ebf",
  1703 => x"f1c21ecc",
  1704 => x"49bf97f0",
  1705 => x"c187f9ee",
  1706 => x"c049cced",
  1707 => x"f487ffe1",
  1708 => x"1e4f268e",
  1709 => x"48c0edc1",
  1710 => x"e3c250c0",
  1711 => x"ff49bfe0",
  1712 => x"c087c3d5",
  1713 => x"1e4f2648",
  1714 => x"cdc71e73",
  1715 => x"ccf3c287",
  1716 => x"ff50c048",
  1717 => x"ffc348d4",
  1718 => x"d0cac178",
  1719 => x"c6d7fe49",
  1720 => x"dbe2fe87",
  1721 => x"02987087",
  1722 => x"ebfe87cd",
  1723 => x"987087f9",
  1724 => x"c187c402",
  1725 => x"c087c24a",
  1726 => x"029a724a",
  1727 => x"cac187c8",
  1728 => x"d6fe49dc",
  1729 => x"f3c287e1",
  1730 => x"78c048c0",
  1731 => x"48f0f1c2",
  1732 => x"fd4950c0",
  1733 => x"dafe87fc",
  1734 => x"9b4b7087",
  1735 => x"c187cf02",
  1736 => x"c75be8ee",
  1737 => x"87f8de49",
  1738 => x"e0c049c1",
  1739 => x"f2c287d3",
  1740 => x"d9e1c087",
  1741 => x"f8efc087",
  1742 => x"87f5ff87",
  1743 => x"4f264b26",
  1744 => x"00000000",
  1745 => x"00000000",
  1746 => x"00000001",
  1747 => x"000011da",
  1748 => x"00002cd8",
  1749 => x"b4000000",
  1750 => x"000011da",
  1751 => x"00002cf6",
  1752 => x"b4000000",
  1753 => x"000011da",
  1754 => x"00002d14",
  1755 => x"b4000000",
  1756 => x"000011da",
  1757 => x"00002d32",
  1758 => x"b4000000",
  1759 => x"000011da",
  1760 => x"00002d50",
  1761 => x"b4000000",
  1762 => x"000011da",
  1763 => x"00002d6e",
  1764 => x"b4000000",
  1765 => x"000011da",
  1766 => x"00002d8c",
  1767 => x"b4000000",
  1768 => x"00001530",
  1769 => x"00000000",
  1770 => x"b4000000",
  1771 => x"000012d4",
  1772 => x"00000000",
  1773 => x"b4000000",
  1774 => x"000012a0",
  1775 => x"db86fc1e",
  1776 => x"fc7e7087",
  1777 => x"1e4f268e",
  1778 => x"c048f0fe",
  1779 => x"7909cd78",
  1780 => x"1e4f2609",
  1781 => x"49fceec1",
  1782 => x"4f2687ed",
  1783 => x"bff0fe1e",
  1784 => x"1e4f2648",
  1785 => x"c148f0fe",
  1786 => x"1e4f2678",
  1787 => x"c048f0fe",
  1788 => x"1e4f2678",
  1789 => x"52c04a71",
  1790 => x"0e4f2651",
  1791 => x"5d5c5b5e",
  1792 => x"7186f40e",
  1793 => x"7e6d974d",
  1794 => x"974ca5c1",
  1795 => x"a6c8486c",
  1796 => x"c4486e58",
  1797 => x"c505a866",
  1798 => x"c048ff87",
  1799 => x"caff87e6",
  1800 => x"49a5c287",
  1801 => x"714b6c97",
  1802 => x"6b974ba3",
  1803 => x"7e6c974b",
  1804 => x"80c1486e",
  1805 => x"c758a6c8",
  1806 => x"58a6cc98",
  1807 => x"fe7c9770",
  1808 => x"487387e1",
  1809 => x"4d268ef4",
  1810 => x"4b264c26",
  1811 => x"731e4f26",
  1812 => x"fe86f41e",
  1813 => x"bfe087d5",
  1814 => x"e0c0494b",
  1815 => x"c00299c0",
  1816 => x"4a7387ea",
  1817 => x"c29affc3",
  1818 => x"bf97c0f7",
  1819 => x"c2f7c249",
  1820 => x"c2517281",
  1821 => x"bf97c0f7",
  1822 => x"c1486e7e",
  1823 => x"58a6c880",
  1824 => x"a6cc98c7",
  1825 => x"c0f7c258",
  1826 => x"5066c848",
  1827 => x"7087cdfd",
  1828 => x"87cffd7e",
  1829 => x"4b268ef4",
  1830 => x"c21e4f26",
  1831 => x"fd49c0f7",
  1832 => x"f1c187d1",
  1833 => x"defc49ce",
  1834 => x"87e8c487",
  1835 => x"5e0e4f26",
  1836 => x"0e5d5c5b",
  1837 => x"7e7186fc",
  1838 => x"c24dd4ff",
  1839 => x"fc49c0f7",
  1840 => x"4b7087f9",
  1841 => x"04abb7c0",
  1842 => x"c387f5c2",
  1843 => x"c905abf0",
  1844 => x"ccf6c187",
  1845 => x"c278c148",
  1846 => x"e0c387d6",
  1847 => x"87c905ab",
  1848 => x"48d0f6c1",
  1849 => x"c7c278c1",
  1850 => x"d0f6c187",
  1851 => x"87c602bf",
  1852 => x"4ca3c0c2",
  1853 => x"4c7387c2",
  1854 => x"bfccf6c1",
  1855 => x"87e0c002",
  1856 => x"b7c44974",
  1857 => x"f6c19129",
  1858 => x"4a7481d4",
  1859 => x"92c29acf",
  1860 => x"307248c1",
  1861 => x"baff4a70",
  1862 => x"98694872",
  1863 => x"87db7970",
  1864 => x"b7c44974",
  1865 => x"f6c19129",
  1866 => x"4a7481d4",
  1867 => x"92c29acf",
  1868 => x"307248c3",
  1869 => x"69484a70",
  1870 => x"6e7970b0",
  1871 => x"87e4c005",
  1872 => x"c848d0ff",
  1873 => x"7dc578e1",
  1874 => x"bfd0f6c1",
  1875 => x"c387c302",
  1876 => x"f6c17de0",
  1877 => x"c302bfcc",
  1878 => x"7df0c387",
  1879 => x"d0ff7d73",
  1880 => x"78e0c048",
  1881 => x"48d0f6c1",
  1882 => x"f6c178c0",
  1883 => x"78c048cc",
  1884 => x"49c0f7c2",
  1885 => x"7087c4fa",
  1886 => x"abb7c04b",
  1887 => x"87cbfd03",
  1888 => x"8efc48c0",
  1889 => x"4c264d26",
  1890 => x"4f264b26",
  1891 => x"00000000",
  1892 => x"00000000",
  1893 => x"00000000",
  1894 => x"34343434",
  1895 => x"34343434",
  1896 => x"34343434",
  1897 => x"34343434",
  1898 => x"34343434",
  1899 => x"34343434",
  1900 => x"34343434",
  1901 => x"34343434",
  1902 => x"34343434",
  1903 => x"34343434",
  1904 => x"34343434",
  1905 => x"34343434",
  1906 => x"34343434",
  1907 => x"34343434",
  1908 => x"34343434",
  1909 => x"724ac01e",
  1910 => x"c191c449",
  1911 => x"c081d4f6",
  1912 => x"d082c179",
  1913 => x"ee04aab7",
  1914 => x"0e4f2687",
  1915 => x"5d5c5b5e",
  1916 => x"f74d710e",
  1917 => x"4a7587f5",
  1918 => x"922ab7c4",
  1919 => x"82d4f6c1",
  1920 => x"9ccf4c75",
  1921 => x"496a94c2",
  1922 => x"c32b744b",
  1923 => x"7448c29b",
  1924 => x"ff4c7030",
  1925 => x"714874bc",
  1926 => x"f77a7098",
  1927 => x"487387c5",
  1928 => x"4c264d26",
  1929 => x"4f264b26",
  1930 => x"48d0ff1e",
  1931 => x"7178e1c8",
  1932 => x"08d4ff48",
  1933 => x"1e4f2678",
  1934 => x"c848d0ff",
  1935 => x"487178e1",
  1936 => x"7808d4ff",
  1937 => x"ff4866c4",
  1938 => x"267808d4",
  1939 => x"4a711e4f",
  1940 => x"1e4966c4",
  1941 => x"deff4972",
  1942 => x"48d0ff87",
  1943 => x"fc78e0c0",
  1944 => x"1e4f268e",
  1945 => x"4a711e73",
  1946 => x"abb7c24b",
  1947 => x"a387c803",
  1948 => x"ffc34a49",
  1949 => x"ce87c79a",
  1950 => x"c34a49a3",
  1951 => x"66c89aff",
  1952 => x"49721e49",
  1953 => x"fc87c6ff",
  1954 => x"264b268e",
  1955 => x"d0ff1e4f",
  1956 => x"78c9c848",
  1957 => x"d4ff4871",
  1958 => x"4f267808",
  1959 => x"494a711e",
  1960 => x"d0ff87eb",
  1961 => x"2678c848",
  1962 => x"1e731e4f",
  1963 => x"f7c24b71",
  1964 => x"c302bfd8",
  1965 => x"87ebc287",
  1966 => x"c848d0ff",
  1967 => x"487378c9",
  1968 => x"ffb0e0c0",
  1969 => x"c27808d4",
  1970 => x"c048ccf7",
  1971 => x"0266c878",
  1972 => x"ffc387c5",
  1973 => x"c087c249",
  1974 => x"d4f7c249",
  1975 => x"0266cc59",
  1976 => x"d5c587c6",
  1977 => x"87c44ad5",
  1978 => x"4affffcf",
  1979 => x"5ad8f7c2",
  1980 => x"48d8f7c2",
  1981 => x"4b2678c1",
  1982 => x"5e0e4f26",
  1983 => x"0e5d5c5b",
  1984 => x"f7c24d71",
  1985 => x"754bbfd4",
  1986 => x"87cb029d",
  1987 => x"c191c849",
  1988 => x"714ae0fa",
  1989 => x"c187c482",
  1990 => x"c04ae0fe",
  1991 => x"7349124c",
  1992 => x"d0f7c299",
  1993 => x"b87148bf",
  1994 => x"7808d4ff",
  1995 => x"842bb7c1",
  1996 => x"04acb7c8",
  1997 => x"f7c287e7",
  1998 => x"c848bfcc",
  1999 => x"d0f7c280",
  2000 => x"264d2658",
  2001 => x"264b264c",
  2002 => x"1e731e4f",
  2003 => x"4a134b71",
  2004 => x"87cb029a",
  2005 => x"e1fe4972",
  2006 => x"9a4a1387",
  2007 => x"2687f505",
  2008 => x"1e4f264b",
  2009 => x"bfccf7c2",
  2010 => x"ccf7c249",
  2011 => x"78a1c148",
  2012 => x"a9b7c0c4",
  2013 => x"ff87db03",
  2014 => x"f7c248d4",
  2015 => x"c278bfd0",
  2016 => x"49bfccf7",
  2017 => x"48ccf7c2",
  2018 => x"c478a1c1",
  2019 => x"04a9b7c0",
  2020 => x"d0ff87e5",
  2021 => x"c278c848",
  2022 => x"c048d8f7",
  2023 => x"004f2678",
  2024 => x"00000000",
  2025 => x"00000000",
  2026 => x"5f000000",
  2027 => x"0000005f",
  2028 => x"00030300",
  2029 => x"00000303",
  2030 => x"147f7f14",
  2031 => x"00147f7f",
  2032 => x"6b2e2400",
  2033 => x"00123a6b",
  2034 => x"18366a4c",
  2035 => x"0032566c",
  2036 => x"594f7e30",
  2037 => x"40683a77",
  2038 => x"07040000",
  2039 => x"00000003",
  2040 => x"3e1c0000",
  2041 => x"00004163",
  2042 => x"63410000",
  2043 => x"00001c3e",
  2044 => x"1c3e2a08",
  2045 => x"082a3e1c",
  2046 => x"3e080800",
  2047 => x"0008083e",
  2048 => x"e0800000",
  2049 => x"00000060",
  2050 => x"08080800",
  2051 => x"00080808",
  2052 => x"60000000",
  2053 => x"00000060",
  2054 => x"18306040",
  2055 => x"0103060c",
  2056 => x"597f3e00",
  2057 => x"003e7f4d",
  2058 => x"7f060400",
  2059 => x"0000007f",
  2060 => x"71634200",
  2061 => x"00464f59",
  2062 => x"49632200",
  2063 => x"00367f49",
  2064 => x"13161c18",
  2065 => x"00107f7f",
  2066 => x"45672700",
  2067 => x"00397d45",
  2068 => x"4b7e3c00",
  2069 => x"00307949",
  2070 => x"71010100",
  2071 => x"00070f79",
  2072 => x"497f3600",
  2073 => x"00367f49",
  2074 => x"494f0600",
  2075 => x"001e3f69",
  2076 => x"66000000",
  2077 => x"00000066",
  2078 => x"e6800000",
  2079 => x"00000066",
  2080 => x"14080800",
  2081 => x"00222214",
  2082 => x"14141400",
  2083 => x"00141414",
  2084 => x"14222200",
  2085 => x"00080814",
  2086 => x"51030200",
  2087 => x"00060f59",
  2088 => x"5d417f3e",
  2089 => x"001e1f55",
  2090 => x"097f7e00",
  2091 => x"007e7f09",
  2092 => x"497f7f00",
  2093 => x"00367f49",
  2094 => x"633e1c00",
  2095 => x"00414141",
  2096 => x"417f7f00",
  2097 => x"001c3e63",
  2098 => x"497f7f00",
  2099 => x"00414149",
  2100 => x"097f7f00",
  2101 => x"00010109",
  2102 => x"417f3e00",
  2103 => x"007a7b49",
  2104 => x"087f7f00",
  2105 => x"007f7f08",
  2106 => x"7f410000",
  2107 => x"0000417f",
  2108 => x"40602000",
  2109 => x"003f7f40",
  2110 => x"1c087f7f",
  2111 => x"00416336",
  2112 => x"407f7f00",
  2113 => x"00404040",
  2114 => x"0c067f7f",
  2115 => x"007f7f06",
  2116 => x"0c067f7f",
  2117 => x"007f7f18",
  2118 => x"417f3e00",
  2119 => x"003e7f41",
  2120 => x"097f7f00",
  2121 => x"00060f09",
  2122 => x"61417f3e",
  2123 => x"00407e7f",
  2124 => x"097f7f00",
  2125 => x"00667f19",
  2126 => x"4d6f2600",
  2127 => x"00327b59",
  2128 => x"7f010100",
  2129 => x"0001017f",
  2130 => x"407f3f00",
  2131 => x"003f7f40",
  2132 => x"703f0f00",
  2133 => x"000f3f70",
  2134 => x"18307f7f",
  2135 => x"007f7f30",
  2136 => x"1c366341",
  2137 => x"4163361c",
  2138 => x"7c060301",
  2139 => x"0103067c",
  2140 => x"4d597161",
  2141 => x"00414347",
  2142 => x"7f7f0000",
  2143 => x"00004141",
  2144 => x"0c060301",
  2145 => x"40603018",
  2146 => x"41410000",
  2147 => x"00007f7f",
  2148 => x"03060c08",
  2149 => x"00080c06",
  2150 => x"80808080",
  2151 => x"00808080",
  2152 => x"03000000",
  2153 => x"00000407",
  2154 => x"54742000",
  2155 => x"00787c54",
  2156 => x"447f7f00",
  2157 => x"00387c44",
  2158 => x"447c3800",
  2159 => x"00004444",
  2160 => x"447c3800",
  2161 => x"007f7f44",
  2162 => x"547c3800",
  2163 => x"00185c54",
  2164 => x"7f7e0400",
  2165 => x"00000505",
  2166 => x"a4bc1800",
  2167 => x"007cfca4",
  2168 => x"047f7f00",
  2169 => x"00787c04",
  2170 => x"3d000000",
  2171 => x"0000407d",
  2172 => x"80808000",
  2173 => x"00007dfd",
  2174 => x"107f7f00",
  2175 => x"00446c38",
  2176 => x"3f000000",
  2177 => x"0000407f",
  2178 => x"180c7c7c",
  2179 => x"00787c0c",
  2180 => x"047c7c00",
  2181 => x"00787c04",
  2182 => x"447c3800",
  2183 => x"00387c44",
  2184 => x"24fcfc00",
  2185 => x"00183c24",
  2186 => x"243c1800",
  2187 => x"00fcfc24",
  2188 => x"047c7c00",
  2189 => x"00080c04",
  2190 => x"545c4800",
  2191 => x"00207454",
  2192 => x"7f3f0400",
  2193 => x"00004444",
  2194 => x"407c3c00",
  2195 => x"007c7c40",
  2196 => x"603c1c00",
  2197 => x"001c3c60",
  2198 => x"30607c3c",
  2199 => x"003c7c60",
  2200 => x"10386c44",
  2201 => x"00446c38",
  2202 => x"e0bc1c00",
  2203 => x"001c3c60",
  2204 => x"74644400",
  2205 => x"00444c5c",
  2206 => x"3e080800",
  2207 => x"00414177",
  2208 => x"7f000000",
  2209 => x"0000007f",
  2210 => x"77414100",
  2211 => x"0008083e",
  2212 => x"03010102",
  2213 => x"00010202",
  2214 => x"7f7f7f7f",
  2215 => x"007f7f7f",
  2216 => x"1c1c0808",
  2217 => x"7f7f3e3e",
  2218 => x"3e3e7f7f",
  2219 => x"08081c1c",
  2220 => x"7c181000",
  2221 => x"0010187c",
  2222 => x"7c301000",
  2223 => x"0010307c",
  2224 => x"60603010",
  2225 => x"00061e78",
  2226 => x"183c6642",
  2227 => x"0042663c",
  2228 => x"c26a3878",
  2229 => x"00386cc6",
  2230 => x"60000060",
  2231 => x"00600000",
  2232 => x"5c5b5e0e",
  2233 => x"86fc0e5d",
  2234 => x"f7c27e71",
  2235 => x"c04cbfe0",
  2236 => x"c41ec04b",
  2237 => x"c402ab66",
  2238 => x"c24dc087",
  2239 => x"754dc187",
  2240 => x"ee49731e",
  2241 => x"86c887e3",
  2242 => x"ef49e0c0",
  2243 => x"a4c487ec",
  2244 => x"f0496a4a",
  2245 => x"caf187f3",
  2246 => x"c184cc87",
  2247 => x"abb7c883",
  2248 => x"87cdff04",
  2249 => x"4d268efc",
  2250 => x"4b264c26",
  2251 => x"711e4f26",
  2252 => x"e4f7c24a",
  2253 => x"e4f7c25a",
  2254 => x"4978c748",
  2255 => x"2687e1fe",
  2256 => x"1e731e4f",
  2257 => x"0bfc4b71",
  2258 => x"4a730b7b",
  2259 => x"c0c19ac1",
  2260 => x"c7ed49a2",
  2261 => x"d8dac287",
  2262 => x"264b265b",
  2263 => x"4a711e4f",
  2264 => x"721e66c4",
  2265 => x"87fbeb49",
  2266 => x"4f268efc",
  2267 => x"48d4ff1e",
  2268 => x"ff78ffc3",
  2269 => x"e1c048d0",
  2270 => x"48d4ff78",
  2271 => x"487178c1",
  2272 => x"d4ff30c4",
  2273 => x"d0ff7808",
  2274 => x"78e0c048",
  2275 => x"5e0e4f26",
  2276 => x"0e5d5c5b",
  2277 => x"7ec086f4",
  2278 => x"ec48a6c8",
  2279 => x"80fc78bf",
  2280 => x"bfe0f7c2",
  2281 => x"e8f7c278",
  2282 => x"bfe84cbf",
  2283 => x"d4dac24d",
  2284 => x"f9e349bf",
  2285 => x"e849c787",
  2286 => x"497087f1",
  2287 => x"d00599c2",
  2288 => x"ccdac287",
  2289 => x"b9ff49bf",
  2290 => x"c19966c8",
  2291 => x"f9c10299",
  2292 => x"49e8cf87",
  2293 => x"7087c1cb",
  2294 => x"e849c74b",
  2295 => x"987087cd",
  2296 => x"c887c905",
  2297 => x"99c14966",
  2298 => x"87fec002",
  2299 => x"ec48a6c8",
  2300 => x"f9e278bf",
  2301 => x"ca497387",
  2302 => x"987087ea",
  2303 => x"c287d702",
  2304 => x"49bfc8da",
  2305 => x"dac2b9c1",
  2306 => x"fd7159cc",
  2307 => x"e8cf87de",
  2308 => x"87c4ca49",
  2309 => x"49c74b70",
  2310 => x"7087d0e7",
  2311 => x"cbff0598",
  2312 => x"4966c887",
  2313 => x"ff0599c1",
  2314 => x"dac287c2",
  2315 => x"c14abfd4",
  2316 => x"d8dac2ba",
  2317 => x"7a0afc5a",
  2318 => x"c19ac10a",
  2319 => x"e949a2c0",
  2320 => x"dac187da",
  2321 => x"87e3e649",
  2322 => x"dac27ec1",
  2323 => x"66c848cc",
  2324 => x"d4dac278",
  2325 => x"e9c005bf",
  2326 => x"c3497587",
  2327 => x"1e7199ff",
  2328 => x"f8fb49c0",
  2329 => x"c8497587",
  2330 => x"1e7129b7",
  2331 => x"ecfb49c1",
  2332 => x"c386c887",
  2333 => x"f2e549fd",
  2334 => x"49fac387",
  2335 => x"c787ece5",
  2336 => x"497587f5",
  2337 => x"c899ffc3",
  2338 => x"b5712db7",
  2339 => x"c0029d75",
  2340 => x"a6c887e4",
  2341 => x"bfc8ff48",
  2342 => x"4966c878",
  2343 => x"bfd0dac2",
  2344 => x"a9e0c289",
  2345 => x"87c4c003",
  2346 => x"87d04dc0",
  2347 => x"48d0dac2",
  2348 => x"c07866c8",
  2349 => x"dac287c6",
  2350 => x"78c048d0",
  2351 => x"99c84975",
  2352 => x"87cec005",
  2353 => x"e449f5c3",
  2354 => x"497087e1",
  2355 => x"c00299c2",
  2356 => x"f7c287e7",
  2357 => x"c002bfe4",
  2358 => x"c14887ca",
  2359 => x"e8f7c288",
  2360 => x"87d3c058",
  2361 => x"c14866c4",
  2362 => x"7e7080e0",
  2363 => x"c002bf6e",
  2364 => x"ff4b87c5",
  2365 => x"c10f7349",
  2366 => x"c449757e",
  2367 => x"cec00599",
  2368 => x"49f2c387",
  2369 => x"7087e4e3",
  2370 => x"0299c249",
  2371 => x"c287ebc0",
  2372 => x"7ebfe4f7",
  2373 => x"b7c7486e",
  2374 => x"cbc003a8",
  2375 => x"c1486e87",
  2376 => x"e8f7c280",
  2377 => x"87d0c058",
  2378 => x"c14a66c4",
  2379 => x"026a82e0",
  2380 => x"4b87c5c0",
  2381 => x"0f7349fe",
  2382 => x"fdc37ec1",
  2383 => x"87ebe249",
  2384 => x"99c24970",
  2385 => x"87e6c002",
  2386 => x"bfe4f7c2",
  2387 => x"87c9c002",
  2388 => x"48e4f7c2",
  2389 => x"d3c078c0",
  2390 => x"4866c487",
  2391 => x"7080e0c1",
  2392 => x"02bf6e7e",
  2393 => x"4b87c5c0",
  2394 => x"0f7349fd",
  2395 => x"fac37ec1",
  2396 => x"87f7e149",
  2397 => x"99c24970",
  2398 => x"87eac002",
  2399 => x"bfe4f7c2",
  2400 => x"a8b7c748",
  2401 => x"87c9c003",
  2402 => x"48e4f7c2",
  2403 => x"d3c078c7",
  2404 => x"4866c487",
  2405 => x"7080e0c1",
  2406 => x"02bf6e7e",
  2407 => x"4b87c5c0",
  2408 => x"0f7349fc",
  2409 => x"48757ec1",
  2410 => x"cc98f0c3",
  2411 => x"987058a6",
  2412 => x"87cec005",
  2413 => x"e049dac1",
  2414 => x"497087f1",
  2415 => x"c10299c2",
  2416 => x"e8cf87f9",
  2417 => x"87d0c349",
  2418 => x"f7c24b70",
  2419 => x"50c048dc",
  2420 => x"97dcf7c2",
  2421 => x"d2c105bf",
  2422 => x"0566c887",
  2423 => x"c187ccc0",
  2424 => x"c6e049da",
  2425 => x"02987087",
  2426 => x"e887c0c1",
  2427 => x"c3494dbf",
  2428 => x"b7c899ff",
  2429 => x"ffb5712d",
  2430 => x"7387f3da",
  2431 => x"87e4c249",
  2432 => x"c0029870",
  2433 => x"f7c287c6",
  2434 => x"50c148dc",
  2435 => x"97dcf7c2",
  2436 => x"d6c005bf",
  2437 => x"c3497587",
  2438 => x"ff0599f0",
  2439 => x"dac187cd",
  2440 => x"c6dfff49",
  2441 => x"05987087",
  2442 => x"c287c0ff",
  2443 => x"49bfe4f7",
  2444 => x"c493cc4b",
  2445 => x"4b6b8366",
  2446 => x"740f7371",
  2447 => x"e9c0029c",
  2448 => x"c0026c87",
  2449 => x"496c87e4",
  2450 => x"87dfdeff",
  2451 => x"99c14970",
  2452 => x"87cbc002",
  2453 => x"c24ba4c4",
  2454 => x"49bfe4f7",
  2455 => x"c80f4b6b",
  2456 => x"c5c00284",
  2457 => x"ff056c87",
  2458 => x"026e87dc",
  2459 => x"c287c8c0",
  2460 => x"49bfe4f7",
  2461 => x"f487e9f1",
  2462 => x"264d268e",
  2463 => x"264b264c",
  2464 => x"0000004f",
  2465 => x"00000010",
  2466 => x"00000000",
  2467 => x"00000000",
  2468 => x"00000000",
  2469 => x"00000000",
  2470 => x"ff4a711e",
  2471 => x"7249bfc8",
  2472 => x"4f2648a1",
  2473 => x"bfc8ff1e",
  2474 => x"c0c0fe89",
  2475 => x"a9c0c0c0",
  2476 => x"c087c401",
  2477 => x"c187c24a",
  2478 => x"2648724a",
  2479 => x"5b5e0e4f",
  2480 => x"710e5d5c",
  2481 => x"4cd4ff4b",
  2482 => x"c04866d0",
  2483 => x"ff49d678",
  2484 => x"c387d5dd",
  2485 => x"496c7cff",
  2486 => x"7199ffc3",
  2487 => x"f0c3494d",
  2488 => x"a9e0c199",
  2489 => x"c387cb05",
  2490 => x"486c7cff",
  2491 => x"66d098c3",
  2492 => x"ffc37808",
  2493 => x"494a6c7c",
  2494 => x"ffc331c8",
  2495 => x"714a6c7c",
  2496 => x"c84972b2",
  2497 => x"7cffc331",
  2498 => x"b2714a6c",
  2499 => x"31c84972",
  2500 => x"6c7cffc3",
  2501 => x"ffb2714a",
  2502 => x"e0c048d0",
  2503 => x"029b7378",
  2504 => x"7b7287c2",
  2505 => x"4d264875",
  2506 => x"4b264c26",
  2507 => x"261e4f26",
  2508 => x"5b5e0e4f",
  2509 => x"86f80e5c",
  2510 => x"a6c81e76",
  2511 => x"87fdfd49",
  2512 => x"4b7086c4",
  2513 => x"a8c4486e",
  2514 => x"87fbc203",
  2515 => x"f0c34a73",
  2516 => x"aad0c19a",
  2517 => x"c187c702",
  2518 => x"c205aae0",
  2519 => x"497387e9",
  2520 => x"c30299c8",
  2521 => x"87c6ff87",
  2522 => x"9cc34c73",
  2523 => x"c105acc2",
  2524 => x"66c487c4",
  2525 => x"7131c949",
  2526 => x"4a66c41e",
  2527 => x"c292ccc1",
  2528 => x"7249ecf7",
  2529 => x"c1cdfe81",
  2530 => x"ff49d887",
  2531 => x"c887d9da",
  2532 => x"e4c21ec0",
  2533 => x"e6fd49e4",
  2534 => x"d0ff87d9",
  2535 => x"78e0c048",
  2536 => x"1ee4e4c2",
  2537 => x"c14a66cc",
  2538 => x"f7c292cc",
  2539 => x"817249ec",
  2540 => x"87d7cbfe",
  2541 => x"acc186cc",
  2542 => x"87cbc105",
  2543 => x"fd49eec0",
  2544 => x"c487c9e3",
  2545 => x"31c94966",
  2546 => x"66c41e71",
  2547 => x"92ccc14a",
  2548 => x"49ecf7c2",
  2549 => x"cbfe8172",
  2550 => x"e4c287f0",
  2551 => x"66c81ee4",
  2552 => x"92ccc14a",
  2553 => x"49ecf7c2",
  2554 => x"c9fe8172",
  2555 => x"49d787de",
  2556 => x"87f4d8ff",
  2557 => x"c21ec0c8",
  2558 => x"fd49e4e4",
  2559 => x"cc87d1e4",
  2560 => x"48d0ff86",
  2561 => x"f878e0c0",
  2562 => x"264c268e",
  2563 => x"1e4f264b",
  2564 => x"b7c44a71",
  2565 => x"87ce03aa",
  2566 => x"ccc14972",
  2567 => x"ecf7c291",
  2568 => x"81c8c181",
  2569 => x"4f2679c0",
  2570 => x"5c5b5e0e",
  2571 => x"86fc0e5d",
  2572 => x"d4ff4a71",
  2573 => x"d44cc04b",
  2574 => x"b7c34d66",
  2575 => x"c2c201ad",
  2576 => x"029a7287",
  2577 => x"1e87ecc0",
  2578 => x"ccc14975",
  2579 => x"ecf7c291",
  2580 => x"c8807148",
  2581 => x"66c458a6",
  2582 => x"fbc2fe49",
  2583 => x"7086c487",
  2584 => x"87d40298",
  2585 => x"c8c1496e",
  2586 => x"6e79c181",
  2587 => x"6981c849",
  2588 => x"7587c54c",
  2589 => x"87d7fe49",
  2590 => x"c848d0ff",
  2591 => x"7bdd78e1",
  2592 => x"ffc34874",
  2593 => x"747b7098",
  2594 => x"29b7c849",
  2595 => x"ffc34871",
  2596 => x"747b7098",
  2597 => x"29b7d049",
  2598 => x"ffc34871",
  2599 => x"747b7098",
  2600 => x"28b7d848",
  2601 => x"7bc07b70",
  2602 => x"7b7b7b7b",
  2603 => x"7b7b7b7b",
  2604 => x"ff7b7b7b",
  2605 => x"e0c048d0",
  2606 => x"dc1e7578",
  2607 => x"ccd6ff49",
  2608 => x"fc86c487",
  2609 => x"264d268e",
  2610 => x"264b264c",
  2611 => x"0000004f",
  2612 => x"ffffffff",
  2613 => x"ffffffff",
  2614 => x"ffffffff",
  2615 => x"ffffffff",
  2616 => x"000028e4",
  2617 => x"33495653",
  2618 => x"20203832",
  2619 => x"004d4f52",
  2620 => x"00001bd3",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
