
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"dc",x"fc",x"c2",x"87"),
    12 => (x"48",x"c0",x"c8",x"4e"),
    13 => (x"d5",x"c1",x"28",x"c2"),
    14 => (x"ea",x"d6",x"e5",x"ea"),
    15 => (x"c1",x"46",x"71",x"49"),
    16 => (x"87",x"f9",x"01",x"88"),
    17 => (x"49",x"dc",x"fc",x"c2"),
    18 => (x"48",x"f4",x"e3",x"c2"),
    19 => (x"03",x"89",x"d0",x"89"),
    20 => (x"40",x"40",x"40",x"c0"),
    21 => (x"d0",x"87",x"f6",x"40"),
    22 => (x"50",x"c0",x"05",x"81"),
    23 => (x"f9",x"05",x"89",x"c1"),
    24 => (x"f4",x"e3",x"c2",x"87"),
    25 => (x"f0",x"e3",x"c2",x"4d"),
    26 => (x"02",x"ad",x"74",x"4c"),
    27 => (x"0f",x"24",x"87",x"c4"),
    28 => (x"e9",x"c1",x"87",x"f7"),
    29 => (x"e3",x"c2",x"87",x"d1"),
    30 => (x"e3",x"c2",x"4d",x"f4"),
    31 => (x"ad",x"74",x"4c",x"f4"),
    32 => (x"c4",x"87",x"c6",x"02"),
    33 => (x"f5",x"0f",x"6c",x"8c"),
    34 => (x"87",x"fd",x"00",x"87"),
    35 => (x"71",x"86",x"fc",x"1e"),
    36 => (x"49",x"c0",x"ff",x"4a"),
    37 => (x"c0",x"c4",x"48",x"69"),
    38 => (x"48",x"7e",x"70",x"98"),
    39 => (x"87",x"f4",x"02",x"98"),
    40 => (x"fc",x"48",x"79",x"72"),
    41 => (x"0e",x"4f",x"26",x"8e"),
    42 => (x"0e",x"5c",x"5b",x"5e"),
    43 => (x"4c",x"c0",x"4b",x"71"),
    44 => (x"02",x"9a",x"4a",x"13"),
    45 => (x"49",x"72",x"87",x"cd"),
    46 => (x"c1",x"87",x"d1",x"ff"),
    47 => (x"9a",x"4a",x"13",x"84"),
    48 => (x"74",x"87",x"f3",x"05"),
    49 => (x"26",x"4c",x"26",x"48"),
    50 => (x"1e",x"4f",x"26",x"4b"),
    51 => (x"1e",x"73",x"1e",x"72"),
    52 => (x"02",x"11",x"48",x"12"),
    53 => (x"c3",x"4b",x"87",x"ca"),
    54 => (x"73",x"9b",x"98",x"df"),
    55 => (x"87",x"f0",x"02",x"88"),
    56 => (x"4a",x"26",x"4b",x"26"),
    57 => (x"73",x"1e",x"4f",x"26"),
    58 => (x"c1",x"1e",x"72",x"1e"),
    59 => (x"87",x"ca",x"04",x"8b"),
    60 => (x"02",x"11",x"48",x"12"),
    61 => (x"02",x"88",x"87",x"c4"),
    62 => (x"4a",x"26",x"87",x"f1"),
    63 => (x"4f",x"26",x"4b",x"26"),
    64 => (x"81",x"48",x"73",x"1e"),
    65 => (x"c5",x"02",x"a9",x"73"),
    66 => (x"05",x"53",x"12",x"87"),
    67 => (x"4f",x"26",x"87",x"f6"),
    68 => (x"71",x"1e",x"73",x"1e"),
    69 => (x"4b",x"66",x"c8",x"4a"),
    70 => (x"71",x"8b",x"c1",x"49"),
    71 => (x"87",x"cf",x"02",x"99"),
    72 => (x"d4",x"ff",x"48",x"12"),
    73 => (x"49",x"73",x"78",x"08"),
    74 => (x"99",x"71",x"8b",x"c1"),
    75 => (x"26",x"87",x"f1",x"05"),
    76 => (x"0e",x"4f",x"26",x"4b"),
    77 => (x"0e",x"5c",x"5b",x"5e"),
    78 => (x"d4",x"ff",x"4a",x"71"),
    79 => (x"4b",x"66",x"cc",x"4c"),
    80 => (x"71",x"8b",x"c1",x"49"),
    81 => (x"87",x"ce",x"02",x"99"),
    82 => (x"6c",x"7c",x"ff",x"c3"),
    83 => (x"c1",x"49",x"73",x"52"),
    84 => (x"05",x"99",x"71",x"8b"),
    85 => (x"4c",x"26",x"87",x"f2"),
    86 => (x"4f",x"26",x"4b",x"26"),
    87 => (x"ff",x"1e",x"73",x"1e"),
    88 => (x"ff",x"c3",x"4b",x"d4"),
    89 => (x"c3",x"4a",x"6b",x"7b"),
    90 => (x"49",x"6b",x"7b",x"ff"),
    91 => (x"b1",x"72",x"32",x"c8"),
    92 => (x"6b",x"7b",x"ff",x"c3"),
    93 => (x"71",x"31",x"c8",x"4a"),
    94 => (x"7b",x"ff",x"c3",x"b2"),
    95 => (x"32",x"c8",x"49",x"6b"),
    96 => (x"48",x"71",x"b1",x"72"),
    97 => (x"4f",x"26",x"4b",x"26"),
    98 => (x"5c",x"5b",x"5e",x"0e"),
    99 => (x"4d",x"71",x"0e",x"5d"),
   100 => (x"75",x"4c",x"d4",x"ff"),
   101 => (x"98",x"ff",x"c3",x"48"),
   102 => (x"e3",x"c2",x"7c",x"70"),
   103 => (x"c8",x"05",x"bf",x"f4"),
   104 => (x"48",x"66",x"d0",x"87"),
   105 => (x"a6",x"d4",x"30",x"c9"),
   106 => (x"49",x"66",x"d0",x"58"),
   107 => (x"48",x"71",x"29",x"d8"),
   108 => (x"70",x"98",x"ff",x"c3"),
   109 => (x"49",x"66",x"d0",x"7c"),
   110 => (x"48",x"71",x"29",x"d0"),
   111 => (x"70",x"98",x"ff",x"c3"),
   112 => (x"49",x"66",x"d0",x"7c"),
   113 => (x"48",x"71",x"29",x"c8"),
   114 => (x"70",x"98",x"ff",x"c3"),
   115 => (x"48",x"66",x"d0",x"7c"),
   116 => (x"70",x"98",x"ff",x"c3"),
   117 => (x"d0",x"49",x"75",x"7c"),
   118 => (x"c3",x"48",x"71",x"29"),
   119 => (x"7c",x"70",x"98",x"ff"),
   120 => (x"f0",x"c9",x"4b",x"6c"),
   121 => (x"ff",x"c3",x"4a",x"ff"),
   122 => (x"87",x"cf",x"05",x"ab"),
   123 => (x"6c",x"7c",x"71",x"49"),
   124 => (x"02",x"8a",x"c1",x"4b"),
   125 => (x"ab",x"71",x"87",x"c5"),
   126 => (x"73",x"87",x"f2",x"02"),
   127 => (x"26",x"4d",x"26",x"48"),
   128 => (x"26",x"4b",x"26",x"4c"),
   129 => (x"49",x"c0",x"1e",x"4f"),
   130 => (x"c3",x"48",x"d4",x"ff"),
   131 => (x"81",x"c1",x"78",x"ff"),
   132 => (x"a9",x"b7",x"c8",x"c3"),
   133 => (x"26",x"87",x"f1",x"04"),
   134 => (x"5b",x"5e",x"0e",x"4f"),
   135 => (x"c0",x"0e",x"5d",x"5c"),
   136 => (x"f7",x"c1",x"f0",x"ff"),
   137 => (x"c0",x"c0",x"c1",x"4d"),
   138 => (x"4b",x"c0",x"c0",x"c0"),
   139 => (x"c4",x"87",x"d6",x"ff"),
   140 => (x"c0",x"4c",x"df",x"f8"),
   141 => (x"fd",x"49",x"75",x"1e"),
   142 => (x"86",x"c4",x"87",x"ce"),
   143 => (x"c0",x"05",x"a8",x"c1"),
   144 => (x"d4",x"ff",x"87",x"e5"),
   145 => (x"78",x"ff",x"c3",x"48"),
   146 => (x"e1",x"c0",x"1e",x"73"),
   147 => (x"49",x"e9",x"c1",x"f0"),
   148 => (x"c4",x"87",x"f5",x"fc"),
   149 => (x"05",x"98",x"70",x"86"),
   150 => (x"d4",x"ff",x"87",x"ca"),
   151 => (x"78",x"ff",x"c3",x"48"),
   152 => (x"87",x"cb",x"48",x"c1"),
   153 => (x"c1",x"87",x"de",x"fe"),
   154 => (x"c6",x"ff",x"05",x"8c"),
   155 => (x"26",x"48",x"c0",x"87"),
   156 => (x"26",x"4c",x"26",x"4d"),
   157 => (x"0e",x"4f",x"26",x"4b"),
   158 => (x"0e",x"5c",x"5b",x"5e"),
   159 => (x"c1",x"f0",x"ff",x"c0"),
   160 => (x"d4",x"ff",x"4c",x"c1"),
   161 => (x"78",x"ff",x"c3",x"48"),
   162 => (x"f8",x"49",x"fc",x"ca"),
   163 => (x"4b",x"d3",x"87",x"d9"),
   164 => (x"49",x"74",x"1e",x"c0"),
   165 => (x"c4",x"87",x"f1",x"fb"),
   166 => (x"05",x"98",x"70",x"86"),
   167 => (x"d4",x"ff",x"87",x"ca"),
   168 => (x"78",x"ff",x"c3",x"48"),
   169 => (x"87",x"cb",x"48",x"c1"),
   170 => (x"c1",x"87",x"da",x"fd"),
   171 => (x"df",x"ff",x"05",x"8b"),
   172 => (x"26",x"48",x"c0",x"87"),
   173 => (x"26",x"4b",x"26",x"4c"),
   174 => (x"00",x"00",x"00",x"4f"),
   175 => (x"00",x"44",x"4d",x"43"),
   176 => (x"43",x"48",x"44",x"53"),
   177 => (x"69",x"61",x"66",x"20"),
   178 => (x"00",x"0a",x"21",x"6c"),
   179 => (x"52",x"52",x"45",x"49"),
   180 => (x"00",x"00",x"00",x"00"),
   181 => (x"00",x"49",x"50",x"53"),
   182 => (x"74",x"69",x"72",x"57"),
   183 => (x"61",x"66",x"20",x"65"),
   184 => (x"64",x"65",x"6c",x"69"),
   185 => (x"5e",x"0e",x"00",x"0a"),
   186 => (x"0e",x"5d",x"5c",x"5b"),
   187 => (x"ff",x"4d",x"ff",x"c3"),
   188 => (x"d0",x"fc",x"4b",x"d4"),
   189 => (x"1e",x"ea",x"c6",x"87"),
   190 => (x"c1",x"f0",x"e1",x"c0"),
   191 => (x"c7",x"fa",x"49",x"c8"),
   192 => (x"c1",x"86",x"c4",x"87"),
   193 => (x"87",x"c8",x"02",x"a8"),
   194 => (x"c0",x"87",x"ec",x"fd"),
   195 => (x"87",x"e8",x"c1",x"48"),
   196 => (x"70",x"87",x"c9",x"f9"),
   197 => (x"ff",x"ff",x"cf",x"49"),
   198 => (x"a9",x"ea",x"c6",x"99"),
   199 => (x"fd",x"87",x"c8",x"02"),
   200 => (x"48",x"c0",x"87",x"d5"),
   201 => (x"75",x"87",x"d1",x"c1"),
   202 => (x"4c",x"f1",x"c0",x"7b"),
   203 => (x"70",x"87",x"ea",x"fb"),
   204 => (x"ec",x"c0",x"02",x"98"),
   205 => (x"c0",x"1e",x"c0",x"87"),
   206 => (x"fa",x"c1",x"f0",x"ff"),
   207 => (x"87",x"c8",x"f9",x"49"),
   208 => (x"98",x"70",x"86",x"c4"),
   209 => (x"75",x"87",x"da",x"05"),
   210 => (x"75",x"49",x"6b",x"7b"),
   211 => (x"75",x"7b",x"75",x"7b"),
   212 => (x"c1",x"7b",x"75",x"7b"),
   213 => (x"c4",x"02",x"99",x"c0"),
   214 => (x"db",x"48",x"c1",x"87"),
   215 => (x"d7",x"48",x"c0",x"87"),
   216 => (x"05",x"ac",x"c2",x"87"),
   217 => (x"c0",x"cb",x"87",x"ca"),
   218 => (x"87",x"fb",x"f4",x"49"),
   219 => (x"87",x"c8",x"48",x"c0"),
   220 => (x"fe",x"05",x"8c",x"c1"),
   221 => (x"48",x"c0",x"87",x"f6"),
   222 => (x"4c",x"26",x"4d",x"26"),
   223 => (x"4f",x"26",x"4b",x"26"),
   224 => (x"5c",x"5b",x"5e",x"0e"),
   225 => (x"d0",x"ff",x"0e",x"5d"),
   226 => (x"d0",x"e5",x"c0",x"4d"),
   227 => (x"c2",x"4c",x"c0",x"c1"),
   228 => (x"c1",x"48",x"f4",x"e3"),
   229 => (x"49",x"d4",x"cb",x"78"),
   230 => (x"c7",x"87",x"cc",x"f4"),
   231 => (x"f9",x"7d",x"c2",x"4b"),
   232 => (x"7d",x"c3",x"87",x"e3"),
   233 => (x"49",x"74",x"1e",x"c0"),
   234 => (x"c4",x"87",x"dd",x"f7"),
   235 => (x"05",x"a8",x"c1",x"86"),
   236 => (x"c2",x"4b",x"87",x"c1"),
   237 => (x"87",x"cb",x"05",x"ab"),
   238 => (x"f3",x"49",x"cc",x"cb"),
   239 => (x"48",x"c0",x"87",x"e9"),
   240 => (x"c1",x"87",x"f6",x"c0"),
   241 => (x"d4",x"ff",x"05",x"8b"),
   242 => (x"87",x"da",x"fc",x"87"),
   243 => (x"58",x"f8",x"e3",x"c2"),
   244 => (x"cd",x"05",x"98",x"70"),
   245 => (x"c0",x"1e",x"c1",x"87"),
   246 => (x"d0",x"c1",x"f0",x"ff"),
   247 => (x"87",x"e8",x"f6",x"49"),
   248 => (x"d4",x"ff",x"86",x"c4"),
   249 => (x"78",x"ff",x"c3",x"48"),
   250 => (x"c2",x"87",x"ee",x"c4"),
   251 => (x"c2",x"58",x"fc",x"e3"),
   252 => (x"48",x"d4",x"ff",x"7d"),
   253 => (x"c1",x"78",x"ff",x"c3"),
   254 => (x"26",x"4d",x"26",x"48"),
   255 => (x"26",x"4b",x"26",x"4c"),
   256 => (x"5b",x"5e",x"0e",x"4f"),
   257 => (x"71",x"0e",x"5d",x"5c"),
   258 => (x"4c",x"ff",x"c3",x"4d"),
   259 => (x"74",x"4b",x"d4",x"ff"),
   260 => (x"48",x"d0",x"ff",x"7b"),
   261 => (x"74",x"78",x"c3",x"c4"),
   262 => (x"c0",x"1e",x"75",x"7b"),
   263 => (x"d8",x"c1",x"f0",x"ff"),
   264 => (x"87",x"e4",x"f5",x"49"),
   265 => (x"98",x"70",x"86",x"c4"),
   266 => (x"cb",x"87",x"cb",x"02"),
   267 => (x"f6",x"f1",x"49",x"d8"),
   268 => (x"c0",x"48",x"c1",x"87"),
   269 => (x"7b",x"74",x"87",x"ee"),
   270 => (x"c8",x"7b",x"fe",x"c3"),
   271 => (x"66",x"d4",x"1e",x"c0"),
   272 => (x"87",x"cc",x"f3",x"49"),
   273 => (x"7b",x"74",x"86",x"c4"),
   274 => (x"7b",x"74",x"7b",x"74"),
   275 => (x"4a",x"e0",x"da",x"d8"),
   276 => (x"05",x"6b",x"7b",x"74"),
   277 => (x"8a",x"c1",x"87",x"c5"),
   278 => (x"74",x"87",x"f5",x"05"),
   279 => (x"48",x"d0",x"ff",x"7b"),
   280 => (x"48",x"c0",x"78",x"c2"),
   281 => (x"4c",x"26",x"4d",x"26"),
   282 => (x"4f",x"26",x"4b",x"26"),
   283 => (x"5c",x"5b",x"5e",x"0e"),
   284 => (x"86",x"fc",x"0e",x"5d"),
   285 => (x"d4",x"ff",x"4b",x"71"),
   286 => (x"c5",x"7e",x"c0",x"4c"),
   287 => (x"4a",x"df",x"cd",x"ee"),
   288 => (x"6c",x"7c",x"ff",x"c3"),
   289 => (x"a8",x"fe",x"c3",x"48"),
   290 => (x"87",x"f8",x"c0",x"05"),
   291 => (x"9b",x"73",x"4d",x"74"),
   292 => (x"d4",x"87",x"cc",x"02"),
   293 => (x"49",x"73",x"1e",x"66"),
   294 => (x"c4",x"87",x"d8",x"f2"),
   295 => (x"ff",x"87",x"d4",x"86"),
   296 => (x"d1",x"c4",x"48",x"d0"),
   297 => (x"4a",x"66",x"d4",x"78"),
   298 => (x"c1",x"7d",x"ff",x"c3"),
   299 => (x"87",x"f8",x"05",x"8a"),
   300 => (x"c3",x"5a",x"a6",x"d8"),
   301 => (x"73",x"7c",x"7c",x"ff"),
   302 => (x"87",x"c5",x"05",x"9b"),
   303 => (x"d0",x"48",x"d0",x"ff"),
   304 => (x"7e",x"4a",x"c1",x"78"),
   305 => (x"fe",x"05",x"8a",x"c1"),
   306 => (x"48",x"6e",x"87",x"f6"),
   307 => (x"4d",x"26",x"8e",x"fc"),
   308 => (x"4b",x"26",x"4c",x"26"),
   309 => (x"73",x"1e",x"4f",x"26"),
   310 => (x"c0",x"4a",x"71",x"1e"),
   311 => (x"48",x"d4",x"ff",x"4b"),
   312 => (x"ff",x"78",x"ff",x"c3"),
   313 => (x"c3",x"c4",x"48",x"d0"),
   314 => (x"48",x"d4",x"ff",x"78"),
   315 => (x"72",x"78",x"ff",x"c3"),
   316 => (x"f0",x"ff",x"c0",x"1e"),
   317 => (x"f2",x"49",x"d1",x"c1"),
   318 => (x"86",x"c4",x"87",x"ce"),
   319 => (x"d2",x"05",x"98",x"70"),
   320 => (x"1e",x"c0",x"c8",x"87"),
   321 => (x"fd",x"49",x"66",x"cc"),
   322 => (x"86",x"c4",x"87",x"e2"),
   323 => (x"d0",x"ff",x"4b",x"70"),
   324 => (x"73",x"78",x"c2",x"48"),
   325 => (x"26",x"4b",x"26",x"48"),
   326 => (x"5b",x"5e",x"0e",x"4f"),
   327 => (x"c0",x"0e",x"5d",x"5c"),
   328 => (x"f0",x"ff",x"c0",x"1e"),
   329 => (x"f1",x"49",x"c9",x"c1"),
   330 => (x"1e",x"d2",x"87",x"de"),
   331 => (x"49",x"c4",x"e4",x"c2"),
   332 => (x"c8",x"87",x"f9",x"fc"),
   333 => (x"c1",x"4c",x"c0",x"86"),
   334 => (x"ac",x"b7",x"d2",x"84"),
   335 => (x"c2",x"87",x"f8",x"04"),
   336 => (x"bf",x"97",x"c4",x"e4"),
   337 => (x"99",x"c0",x"c3",x"49"),
   338 => (x"05",x"a9",x"c0",x"c1"),
   339 => (x"c2",x"87",x"e7",x"c0"),
   340 => (x"bf",x"97",x"cb",x"e4"),
   341 => (x"c2",x"31",x"d0",x"49"),
   342 => (x"bf",x"97",x"cc",x"e4"),
   343 => (x"72",x"32",x"c8",x"4a"),
   344 => (x"cd",x"e4",x"c2",x"b1"),
   345 => (x"b1",x"4a",x"bf",x"97"),
   346 => (x"ff",x"cf",x"4c",x"71"),
   347 => (x"c1",x"9c",x"ff",x"ff"),
   348 => (x"c1",x"34",x"ca",x"84"),
   349 => (x"e4",x"c2",x"87",x"e7"),
   350 => (x"49",x"bf",x"97",x"cd"),
   351 => (x"99",x"c6",x"31",x"c1"),
   352 => (x"97",x"ce",x"e4",x"c2"),
   353 => (x"b7",x"c7",x"4a",x"bf"),
   354 => (x"c2",x"b1",x"72",x"2a"),
   355 => (x"bf",x"97",x"c9",x"e4"),
   356 => (x"9d",x"cf",x"4d",x"4a"),
   357 => (x"97",x"ca",x"e4",x"c2"),
   358 => (x"9a",x"c3",x"4a",x"bf"),
   359 => (x"e4",x"c2",x"32",x"ca"),
   360 => (x"4b",x"bf",x"97",x"cb"),
   361 => (x"b2",x"73",x"33",x"c2"),
   362 => (x"97",x"cc",x"e4",x"c2"),
   363 => (x"c0",x"c3",x"4b",x"bf"),
   364 => (x"2b",x"b7",x"c6",x"9b"),
   365 => (x"81",x"c2",x"b2",x"73"),
   366 => (x"30",x"71",x"48",x"c1"),
   367 => (x"48",x"c1",x"49",x"70"),
   368 => (x"4d",x"70",x"30",x"75"),
   369 => (x"84",x"c1",x"4c",x"72"),
   370 => (x"c0",x"c8",x"94",x"71"),
   371 => (x"cc",x"06",x"ad",x"b7"),
   372 => (x"b7",x"34",x"c1",x"87"),
   373 => (x"b7",x"c0",x"c8",x"2d"),
   374 => (x"f4",x"ff",x"01",x"ad"),
   375 => (x"26",x"48",x"74",x"87"),
   376 => (x"26",x"4c",x"26",x"4d"),
   377 => (x"0e",x"4f",x"26",x"4b"),
   378 => (x"5d",x"5c",x"5b",x"5e"),
   379 => (x"c2",x"86",x"fc",x"0e"),
   380 => (x"c0",x"48",x"ec",x"ec"),
   381 => (x"e4",x"e4",x"c2",x"78"),
   382 => (x"fb",x"49",x"c0",x"1e"),
   383 => (x"86",x"c4",x"87",x"d8"),
   384 => (x"c5",x"05",x"98",x"70"),
   385 => (x"c9",x"48",x"c0",x"87"),
   386 => (x"4d",x"c0",x"87",x"d4"),
   387 => (x"48",x"e8",x"f1",x"c2"),
   388 => (x"e5",x"c2",x"78",x"c1"),
   389 => (x"e1",x"c0",x"4a",x"da"),
   390 => (x"4b",x"c8",x"49",x"f4"),
   391 => (x"70",x"87",x"c7",x"eb"),
   392 => (x"87",x"c6",x"05",x"98"),
   393 => (x"48",x"e8",x"f1",x"c2"),
   394 => (x"e5",x"c2",x"78",x"c0"),
   395 => (x"e2",x"c0",x"4a",x"f6"),
   396 => (x"4b",x"c8",x"49",x"c0"),
   397 => (x"70",x"87",x"ef",x"ea"),
   398 => (x"87",x"c6",x"05",x"98"),
   399 => (x"48",x"e8",x"f1",x"c2"),
   400 => (x"f1",x"c2",x"78",x"c0"),
   401 => (x"c0",x"02",x"bf",x"e8"),
   402 => (x"eb",x"c2",x"87",x"fe"),
   403 => (x"c2",x"4d",x"bf",x"ea"),
   404 => (x"bf",x"9f",x"e2",x"ec"),
   405 => (x"c5",x"48",x"6e",x"7e"),
   406 => (x"05",x"a8",x"ea",x"d6"),
   407 => (x"eb",x"c2",x"87",x"c7"),
   408 => (x"ce",x"4d",x"bf",x"ea"),
   409 => (x"ca",x"48",x"6e",x"87"),
   410 => (x"02",x"a8",x"d5",x"e9"),
   411 => (x"48",x"c0",x"87",x"c5"),
   412 => (x"c2",x"87",x"eb",x"c7"),
   413 => (x"75",x"1e",x"e4",x"e4"),
   414 => (x"87",x"da",x"f9",x"49"),
   415 => (x"98",x"70",x"86",x"c4"),
   416 => (x"c0",x"87",x"c5",x"05"),
   417 => (x"87",x"d6",x"c7",x"48"),
   418 => (x"4a",x"f6",x"e5",x"c2"),
   419 => (x"49",x"cc",x"e2",x"c0"),
   420 => (x"d1",x"e9",x"4b",x"c8"),
   421 => (x"05",x"98",x"70",x"87"),
   422 => (x"ec",x"c2",x"87",x"c8"),
   423 => (x"78",x"c1",x"48",x"ec"),
   424 => (x"e5",x"c2",x"87",x"d8"),
   425 => (x"e2",x"c0",x"4a",x"da"),
   426 => (x"4b",x"c8",x"49",x"d8"),
   427 => (x"70",x"87",x"f7",x"e8"),
   428 => (x"c5",x"c0",x"02",x"98"),
   429 => (x"c6",x"48",x"c0",x"87"),
   430 => (x"ec",x"c2",x"87",x"e4"),
   431 => (x"49",x"bf",x"97",x"e2"),
   432 => (x"05",x"a9",x"d5",x"c1"),
   433 => (x"c2",x"87",x"cd",x"c0"),
   434 => (x"bf",x"97",x"e3",x"ec"),
   435 => (x"a9",x"ea",x"c2",x"49"),
   436 => (x"87",x"c5",x"c0",x"02"),
   437 => (x"c5",x"c6",x"48",x"c0"),
   438 => (x"e4",x"e4",x"c2",x"87"),
   439 => (x"6e",x"7e",x"bf",x"97"),
   440 => (x"a8",x"e9",x"c3",x"48"),
   441 => (x"87",x"ce",x"c0",x"02"),
   442 => (x"eb",x"c3",x"48",x"6e"),
   443 => (x"c5",x"c0",x"02",x"a8"),
   444 => (x"c5",x"48",x"c0",x"87"),
   445 => (x"e4",x"c2",x"87",x"e8"),
   446 => (x"49",x"bf",x"97",x"ef"),
   447 => (x"cc",x"c0",x"05",x"99"),
   448 => (x"f0",x"e4",x"c2",x"87"),
   449 => (x"c2",x"49",x"bf",x"97"),
   450 => (x"c5",x"c0",x"02",x"a9"),
   451 => (x"c5",x"48",x"c0",x"87"),
   452 => (x"e4",x"c2",x"87",x"cc"),
   453 => (x"48",x"bf",x"97",x"f1"),
   454 => (x"58",x"e8",x"ec",x"c2"),
   455 => (x"c1",x"48",x"4c",x"70"),
   456 => (x"ec",x"ec",x"c2",x"88"),
   457 => (x"f2",x"e4",x"c2",x"58"),
   458 => (x"75",x"49",x"bf",x"97"),
   459 => (x"f3",x"e4",x"c2",x"81"),
   460 => (x"c8",x"4a",x"bf",x"97"),
   461 => (x"7e",x"a1",x"72",x"32"),
   462 => (x"48",x"c4",x"f1",x"c2"),
   463 => (x"e4",x"c2",x"78",x"6e"),
   464 => (x"48",x"bf",x"97",x"f4"),
   465 => (x"58",x"dc",x"f1",x"c2"),
   466 => (x"bf",x"ec",x"ec",x"c2"),
   467 => (x"87",x"d3",x"c2",x"02"),
   468 => (x"4a",x"f6",x"e5",x"c2"),
   469 => (x"49",x"e8",x"e1",x"c0"),
   470 => (x"c9",x"e6",x"4b",x"c8"),
   471 => (x"02",x"98",x"70",x"87"),
   472 => (x"c0",x"87",x"c5",x"c0"),
   473 => (x"87",x"f6",x"c3",x"48"),
   474 => (x"bf",x"e4",x"ec",x"c2"),
   475 => (x"d8",x"f1",x"c2",x"4c"),
   476 => (x"c9",x"e5",x"c2",x"5c"),
   477 => (x"c8",x"49",x"bf",x"97"),
   478 => (x"c8",x"e5",x"c2",x"31"),
   479 => (x"a1",x"4a",x"bf",x"97"),
   480 => (x"ca",x"e5",x"c2",x"49"),
   481 => (x"d0",x"4a",x"bf",x"97"),
   482 => (x"49",x"a1",x"72",x"32"),
   483 => (x"97",x"cb",x"e5",x"c2"),
   484 => (x"32",x"d8",x"4a",x"bf"),
   485 => (x"c2",x"49",x"a1",x"72"),
   486 => (x"c2",x"59",x"e0",x"f1"),
   487 => (x"91",x"bf",x"d8",x"f1"),
   488 => (x"bf",x"c4",x"f1",x"c2"),
   489 => (x"cc",x"f1",x"c2",x"81"),
   490 => (x"d1",x"e5",x"c2",x"59"),
   491 => (x"c8",x"4a",x"bf",x"97"),
   492 => (x"d0",x"e5",x"c2",x"32"),
   493 => (x"a2",x"4b",x"bf",x"97"),
   494 => (x"d2",x"e5",x"c2",x"4a"),
   495 => (x"d0",x"4b",x"bf",x"97"),
   496 => (x"4a",x"a2",x"73",x"33"),
   497 => (x"97",x"d3",x"e5",x"c2"),
   498 => (x"9b",x"cf",x"4b",x"bf"),
   499 => (x"a2",x"73",x"33",x"d8"),
   500 => (x"d0",x"f1",x"c2",x"4a"),
   501 => (x"74",x"8a",x"c2",x"5a"),
   502 => (x"d0",x"f1",x"c2",x"92"),
   503 => (x"78",x"a1",x"72",x"48"),
   504 => (x"c2",x"87",x"c7",x"c1"),
   505 => (x"bf",x"97",x"f6",x"e4"),
   506 => (x"c2",x"31",x"c8",x"49"),
   507 => (x"bf",x"97",x"f5",x"e4"),
   508 => (x"c5",x"49",x"a1",x"4a"),
   509 => (x"81",x"ff",x"c7",x"31"),
   510 => (x"f1",x"c2",x"29",x"c9"),
   511 => (x"e4",x"c2",x"59",x"d8"),
   512 => (x"4a",x"bf",x"97",x"fb"),
   513 => (x"e4",x"c2",x"32",x"c8"),
   514 => (x"4b",x"bf",x"97",x"fa"),
   515 => (x"f1",x"c2",x"4a",x"a2"),
   516 => (x"f1",x"c2",x"5a",x"e0"),
   517 => (x"6e",x"92",x"bf",x"d8"),
   518 => (x"d4",x"f1",x"c2",x"82"),
   519 => (x"cc",x"f1",x"c2",x"5a"),
   520 => (x"c2",x"78",x"c0",x"48"),
   521 => (x"72",x"48",x"c8",x"f1"),
   522 => (x"f1",x"c2",x"78",x"a1"),
   523 => (x"f1",x"c2",x"48",x"e0"),
   524 => (x"c2",x"78",x"bf",x"cc"),
   525 => (x"c2",x"48",x"e4",x"f1"),
   526 => (x"78",x"bf",x"d0",x"f1"),
   527 => (x"bf",x"ec",x"ec",x"c2"),
   528 => (x"87",x"c9",x"c0",x"02"),
   529 => (x"30",x"c4",x"48",x"74"),
   530 => (x"c9",x"c0",x"7e",x"70"),
   531 => (x"d4",x"f1",x"c2",x"87"),
   532 => (x"30",x"c4",x"48",x"bf"),
   533 => (x"ec",x"c2",x"7e",x"70"),
   534 => (x"78",x"6e",x"48",x"f0"),
   535 => (x"8e",x"fc",x"48",x"c1"),
   536 => (x"4c",x"26",x"4d",x"26"),
   537 => (x"4f",x"26",x"4b",x"26"),
   538 => (x"33",x"54",x"41",x"46"),
   539 => (x"20",x"20",x"20",x"32"),
   540 => (x"00",x"00",x"00",x"00"),
   541 => (x"31",x"54",x"41",x"46"),
   542 => (x"20",x"20",x"20",x"36"),
   543 => (x"00",x"00",x"00",x"00"),
   544 => (x"33",x"54",x"41",x"46"),
   545 => (x"20",x"20",x"20",x"32"),
   546 => (x"00",x"00",x"00",x"00"),
   547 => (x"33",x"54",x"41",x"46"),
   548 => (x"20",x"20",x"20",x"32"),
   549 => (x"00",x"00",x"00",x"00"),
   550 => (x"31",x"54",x"41",x"46"),
   551 => (x"20",x"20",x"20",x"36"),
   552 => (x"5b",x"5e",x"0e",x"00"),
   553 => (x"71",x"0e",x"5d",x"5c"),
   554 => (x"ec",x"ec",x"c2",x"4a"),
   555 => (x"87",x"cb",x"02",x"bf"),
   556 => (x"2b",x"c7",x"4b",x"72"),
   557 => (x"ff",x"c1",x"4d",x"72"),
   558 => (x"72",x"87",x"c9",x"9d"),
   559 => (x"72",x"2b",x"c8",x"4b"),
   560 => (x"9d",x"ff",x"c3",x"4d"),
   561 => (x"bf",x"c4",x"f1",x"c2"),
   562 => (x"ec",x"f9",x"c0",x"83"),
   563 => (x"d9",x"02",x"ab",x"bf"),
   564 => (x"f0",x"f9",x"c0",x"87"),
   565 => (x"e4",x"e4",x"c2",x"5b"),
   566 => (x"ef",x"49",x"73",x"1e"),
   567 => (x"86",x"c4",x"87",x"f8"),
   568 => (x"c5",x"05",x"98",x"70"),
   569 => (x"c0",x"48",x"c0",x"87"),
   570 => (x"ec",x"c2",x"87",x"e6"),
   571 => (x"d2",x"02",x"bf",x"ec"),
   572 => (x"c4",x"49",x"75",x"87"),
   573 => (x"e4",x"e4",x"c2",x"91"),
   574 => (x"cf",x"4c",x"69",x"81"),
   575 => (x"ff",x"ff",x"ff",x"ff"),
   576 => (x"75",x"87",x"cb",x"9c"),
   577 => (x"c2",x"91",x"c2",x"49"),
   578 => (x"9f",x"81",x"e4",x"e4"),
   579 => (x"48",x"74",x"4c",x"69"),
   580 => (x"4c",x"26",x"4d",x"26"),
   581 => (x"4f",x"26",x"4b",x"26"),
   582 => (x"5c",x"5b",x"5e",x"0e"),
   583 => (x"86",x"f4",x"0e",x"5d"),
   584 => (x"c4",x"59",x"a6",x"c8"),
   585 => (x"80",x"c8",x"48",x"66"),
   586 => (x"48",x"6e",x"7e",x"70"),
   587 => (x"c1",x"1e",x"78",x"c0"),
   588 => (x"87",x"fd",x"cc",x"49"),
   589 => (x"4c",x"70",x"86",x"c4"),
   590 => (x"fc",x"c0",x"02",x"9c"),
   591 => (x"f4",x"ec",x"c2",x"87"),
   592 => (x"49",x"66",x"dc",x"4a"),
   593 => (x"87",x"c3",x"de",x"ff"),
   594 => (x"c0",x"02",x"98",x"70"),
   595 => (x"4a",x"74",x"87",x"eb"),
   596 => (x"cb",x"49",x"66",x"dc"),
   597 => (x"cd",x"de",x"ff",x"4b"),
   598 => (x"02",x"98",x"70",x"87"),
   599 => (x"1e",x"c0",x"87",x"db"),
   600 => (x"c4",x"02",x"9c",x"74"),
   601 => (x"c2",x"4d",x"c0",x"87"),
   602 => (x"75",x"4d",x"c1",x"87"),
   603 => (x"87",x"c1",x"cc",x"49"),
   604 => (x"4c",x"70",x"86",x"c4"),
   605 => (x"c4",x"ff",x"05",x"9c"),
   606 => (x"02",x"9c",x"74",x"87"),
   607 => (x"dc",x"87",x"f4",x"c1"),
   608 => (x"48",x"6e",x"49",x"a4"),
   609 => (x"a4",x"da",x"78",x"69"),
   610 => (x"4d",x"66",x"c4",x"49"),
   611 => (x"69",x"9f",x"85",x"c4"),
   612 => (x"ec",x"ec",x"c2",x"7d"),
   613 => (x"87",x"d2",x"02",x"bf"),
   614 => (x"9f",x"49",x"a4",x"d4"),
   615 => (x"ff",x"c0",x"49",x"69"),
   616 => (x"48",x"71",x"99",x"ff"),
   617 => (x"7e",x"70",x"30",x"d0"),
   618 => (x"7e",x"c0",x"87",x"c2"),
   619 => (x"6d",x"48",x"49",x"6e"),
   620 => (x"c4",x"7d",x"70",x"80"),
   621 => (x"78",x"c0",x"48",x"66"),
   622 => (x"cc",x"49",x"66",x"c4"),
   623 => (x"c4",x"79",x"6d",x"81"),
   624 => (x"81",x"d0",x"49",x"66"),
   625 => (x"a6",x"c8",x"79",x"c0"),
   626 => (x"c8",x"78",x"c0",x"48"),
   627 => (x"66",x"c4",x"4c",x"66"),
   628 => (x"74",x"82",x"d4",x"4a"),
   629 => (x"72",x"91",x"c8",x"49"),
   630 => (x"41",x"c0",x"49",x"a1"),
   631 => (x"84",x"c1",x"79",x"6d"),
   632 => (x"04",x"ac",x"b7",x"c6"),
   633 => (x"c4",x"87",x"e7",x"ff"),
   634 => (x"c4",x"c1",x"49",x"66"),
   635 => (x"c1",x"79",x"c0",x"81"),
   636 => (x"c0",x"87",x"c2",x"48"),
   637 => (x"26",x"8e",x"f4",x"48"),
   638 => (x"26",x"4c",x"26",x"4d"),
   639 => (x"0e",x"4f",x"26",x"4b"),
   640 => (x"5d",x"5c",x"5b",x"5e"),
   641 => (x"d0",x"4c",x"71",x"0e"),
   642 => (x"49",x"6c",x"4d",x"66"),
   643 => (x"c2",x"b9",x"75",x"85"),
   644 => (x"4a",x"bf",x"e8",x"ec"),
   645 => (x"99",x"72",x"ba",x"ff"),
   646 => (x"c0",x"02",x"99",x"71"),
   647 => (x"a4",x"c4",x"87",x"e4"),
   648 => (x"f9",x"49",x"6b",x"4b"),
   649 => (x"7b",x"70",x"87",x"fb"),
   650 => (x"bf",x"e4",x"ec",x"c2"),
   651 => (x"71",x"81",x"6c",x"49"),
   652 => (x"c2",x"b9",x"75",x"7c"),
   653 => (x"4a",x"bf",x"e8",x"ec"),
   654 => (x"99",x"72",x"ba",x"ff"),
   655 => (x"ff",x"05",x"99",x"71"),
   656 => (x"7c",x"75",x"87",x"dc"),
   657 => (x"4c",x"26",x"4d",x"26"),
   658 => (x"4f",x"26",x"4b",x"26"),
   659 => (x"71",x"1e",x"73",x"1e"),
   660 => (x"c8",x"f1",x"c2",x"4b"),
   661 => (x"a3",x"c4",x"49",x"bf"),
   662 => (x"c2",x"4a",x"6a",x"4a"),
   663 => (x"e4",x"ec",x"c2",x"8a"),
   664 => (x"a1",x"72",x"92",x"bf"),
   665 => (x"e8",x"ec",x"c2",x"49"),
   666 => (x"9a",x"6b",x"4a",x"bf"),
   667 => (x"c0",x"49",x"a1",x"72"),
   668 => (x"c8",x"59",x"f0",x"f9"),
   669 => (x"e9",x"71",x"1e",x"66"),
   670 => (x"86",x"c4",x"87",x"dc"),
   671 => (x"c4",x"05",x"98",x"70"),
   672 => (x"c2",x"48",x"c0",x"87"),
   673 => (x"26",x"48",x"c1",x"87"),
   674 => (x"1e",x"4f",x"26",x"4b"),
   675 => (x"4b",x"71",x"1e",x"73"),
   676 => (x"bf",x"c8",x"f1",x"c2"),
   677 => (x"4a",x"a3",x"c4",x"49"),
   678 => (x"8a",x"c2",x"4a",x"6a"),
   679 => (x"bf",x"e4",x"ec",x"c2"),
   680 => (x"49",x"a1",x"72",x"92"),
   681 => (x"bf",x"e8",x"ec",x"c2"),
   682 => (x"72",x"9a",x"6b",x"4a"),
   683 => (x"f9",x"c0",x"49",x"a1"),
   684 => (x"66",x"c8",x"59",x"f0"),
   685 => (x"c8",x"e5",x"71",x"1e"),
   686 => (x"70",x"86",x"c4",x"87"),
   687 => (x"87",x"c4",x"05",x"98"),
   688 => (x"87",x"c2",x"48",x"c0"),
   689 => (x"4b",x"26",x"48",x"c1"),
   690 => (x"5e",x"0e",x"4f",x"26"),
   691 => (x"0e",x"5d",x"5c",x"5b"),
   692 => (x"4b",x"71",x"86",x"e4"),
   693 => (x"48",x"66",x"ec",x"c0"),
   694 => (x"a6",x"cc",x"28",x"c9"),
   695 => (x"e8",x"ec",x"c2",x"58"),
   696 => (x"b9",x"ff",x"49",x"bf"),
   697 => (x"66",x"c8",x"48",x"71"),
   698 => (x"58",x"a6",x"d4",x"98"),
   699 => (x"98",x"6b",x"48",x"71"),
   700 => (x"c4",x"58",x"a6",x"d0"),
   701 => (x"a6",x"c4",x"7e",x"a3"),
   702 => (x"78",x"bf",x"6e",x"48"),
   703 => (x"cc",x"48",x"66",x"d0"),
   704 => (x"c6",x"05",x"a8",x"66"),
   705 => (x"7b",x"66",x"c8",x"87"),
   706 => (x"d4",x"87",x"c6",x"c3"),
   707 => (x"ff",x"c1",x"48",x"a6"),
   708 => (x"ff",x"ff",x"ff",x"ff"),
   709 => (x"ff",x"80",x"c4",x"78"),
   710 => (x"d4",x"4a",x"c0",x"78"),
   711 => (x"49",x"72",x"4d",x"a3"),
   712 => (x"a1",x"75",x"91",x"c8"),
   713 => (x"4c",x"66",x"d0",x"49"),
   714 => (x"b7",x"c0",x"8c",x"69"),
   715 => (x"87",x"cd",x"04",x"ac"),
   716 => (x"ac",x"b7",x"66",x"d4"),
   717 => (x"dc",x"87",x"c6",x"03"),
   718 => (x"a6",x"d8",x"5a",x"a6"),
   719 => (x"c6",x"82",x"c1",x"5c"),
   720 => (x"ff",x"04",x"aa",x"b7"),
   721 => (x"66",x"d8",x"87",x"d5"),
   722 => (x"a8",x"b7",x"c0",x"48"),
   723 => (x"d8",x"87",x"d0",x"04"),
   724 => (x"91",x"c8",x"49",x"66"),
   725 => (x"21",x"49",x"a1",x"75"),
   726 => (x"69",x"48",x"6e",x"7b"),
   727 => (x"c0",x"87",x"c9",x"78"),
   728 => (x"49",x"a3",x"cc",x"7b"),
   729 => (x"78",x"69",x"48",x"6e"),
   730 => (x"6b",x"48",x"66",x"c8"),
   731 => (x"58",x"a6",x"cc",x"88"),
   732 => (x"bf",x"e4",x"ec",x"c2"),
   733 => (x"70",x"90",x"c8",x"48"),
   734 => (x"48",x"66",x"c8",x"7e"),
   735 => (x"c9",x"01",x"a8",x"6e"),
   736 => (x"48",x"66",x"c8",x"87"),
   737 => (x"c0",x"03",x"a8",x"6e"),
   738 => (x"c4",x"c1",x"87",x"fd"),
   739 => (x"bf",x"6e",x"7e",x"a3"),
   740 => (x"75",x"91",x"c8",x"49"),
   741 => (x"66",x"cc",x"49",x"a1"),
   742 => (x"49",x"bf",x"6e",x"79"),
   743 => (x"a1",x"75",x"91",x"c8"),
   744 => (x"66",x"81",x"c4",x"49"),
   745 => (x"48",x"a6",x"d0",x"79"),
   746 => (x"d0",x"78",x"bf",x"6e"),
   747 => (x"a8",x"c5",x"48",x"66"),
   748 => (x"c4",x"87",x"c7",x"05"),
   749 => (x"78",x"c0",x"48",x"a6"),
   750 => (x"66",x"d0",x"87",x"c8"),
   751 => (x"c8",x"80",x"c1",x"48"),
   752 => (x"48",x"6e",x"58",x"a6"),
   753 => (x"c8",x"78",x"66",x"c4"),
   754 => (x"49",x"73",x"1e",x"66"),
   755 => (x"c4",x"87",x"f0",x"f8"),
   756 => (x"e4",x"e4",x"c2",x"86"),
   757 => (x"f9",x"49",x"73",x"1e"),
   758 => (x"a3",x"d0",x"87",x"f2"),
   759 => (x"66",x"f0",x"c0",x"49"),
   760 => (x"26",x"8e",x"e0",x"79"),
   761 => (x"26",x"4c",x"26",x"4d"),
   762 => (x"0e",x"4f",x"26",x"4b"),
   763 => (x"0e",x"5c",x"5b",x"5e"),
   764 => (x"4b",x"c0",x"4a",x"71"),
   765 => (x"c0",x"02",x"9a",x"72"),
   766 => (x"a2",x"da",x"87",x"e0"),
   767 => (x"4b",x"69",x"9f",x"49"),
   768 => (x"bf",x"ec",x"ec",x"c2"),
   769 => (x"d4",x"87",x"cf",x"02"),
   770 => (x"69",x"9f",x"49",x"a2"),
   771 => (x"ff",x"c0",x"4c",x"49"),
   772 => (x"34",x"d0",x"9c",x"ff"),
   773 => (x"4c",x"c0",x"87",x"c2"),
   774 => (x"9b",x"73",x"b3",x"74"),
   775 => (x"4a",x"87",x"df",x"02"),
   776 => (x"ec",x"c2",x"8a",x"c2"),
   777 => (x"92",x"49",x"bf",x"e4"),
   778 => (x"bf",x"c8",x"f1",x"c2"),
   779 => (x"c2",x"80",x"72",x"48"),
   780 => (x"71",x"58",x"e8",x"f1"),
   781 => (x"c2",x"30",x"c4",x"48"),
   782 => (x"c0",x"58",x"f4",x"ec"),
   783 => (x"f1",x"c2",x"87",x"e9"),
   784 => (x"c2",x"4b",x"bf",x"cc"),
   785 => (x"c2",x"48",x"e4",x"f1"),
   786 => (x"78",x"bf",x"d0",x"f1"),
   787 => (x"bf",x"ec",x"ec",x"c2"),
   788 => (x"c2",x"87",x"c9",x"02"),
   789 => (x"49",x"bf",x"e4",x"ec"),
   790 => (x"87",x"c7",x"31",x"c4"),
   791 => (x"bf",x"d4",x"f1",x"c2"),
   792 => (x"c2",x"31",x"c4",x"49"),
   793 => (x"c2",x"59",x"f4",x"ec"),
   794 => (x"26",x"5b",x"e4",x"f1"),
   795 => (x"26",x"4b",x"26",x"4c"),
   796 => (x"5b",x"5e",x"0e",x"4f"),
   797 => (x"f0",x"0e",x"5d",x"5c"),
   798 => (x"59",x"a6",x"c8",x"86"),
   799 => (x"ff",x"ff",x"ff",x"cf"),
   800 => (x"7e",x"c0",x"4c",x"f8"),
   801 => (x"d8",x"02",x"66",x"c4"),
   802 => (x"e0",x"e4",x"c2",x"87"),
   803 => (x"c2",x"78",x"c0",x"48"),
   804 => (x"c2",x"48",x"d8",x"e4"),
   805 => (x"78",x"bf",x"e4",x"f1"),
   806 => (x"48",x"dc",x"e4",x"c2"),
   807 => (x"bf",x"e0",x"f1",x"c2"),
   808 => (x"c1",x"ed",x"c2",x"78"),
   809 => (x"c2",x"50",x"c0",x"48"),
   810 => (x"49",x"bf",x"f0",x"ec"),
   811 => (x"bf",x"e0",x"e4",x"c2"),
   812 => (x"03",x"aa",x"71",x"4a"),
   813 => (x"72",x"87",x"cc",x"c4"),
   814 => (x"05",x"99",x"cf",x"49"),
   815 => (x"c0",x"87",x"ea",x"c0"),
   816 => (x"c2",x"48",x"ec",x"f9"),
   817 => (x"78",x"bf",x"d8",x"e4"),
   818 => (x"1e",x"e4",x"e4",x"c2"),
   819 => (x"bf",x"d8",x"e4",x"c2"),
   820 => (x"d8",x"e4",x"c2",x"49"),
   821 => (x"78",x"a1",x"c1",x"48"),
   822 => (x"f9",x"df",x"ff",x"71"),
   823 => (x"c0",x"86",x"c4",x"87"),
   824 => (x"c2",x"48",x"e8",x"f9"),
   825 => (x"cc",x"78",x"e4",x"e4"),
   826 => (x"e8",x"f9",x"c0",x"87"),
   827 => (x"e0",x"c0",x"48",x"bf"),
   828 => (x"ec",x"f9",x"c0",x"80"),
   829 => (x"e0",x"e4",x"c2",x"58"),
   830 => (x"80",x"c1",x"48",x"bf"),
   831 => (x"58",x"e4",x"e4",x"c2"),
   832 => (x"00",x"0e",x"68",x"27"),
   833 => (x"bf",x"97",x"bf",x"00"),
   834 => (x"c2",x"02",x"9d",x"4d"),
   835 => (x"e5",x"c3",x"87",x"e5"),
   836 => (x"de",x"c2",x"02",x"ad"),
   837 => (x"e8",x"f9",x"c0",x"87"),
   838 => (x"a3",x"cb",x"4b",x"bf"),
   839 => (x"cf",x"4c",x"11",x"49"),
   840 => (x"d2",x"c1",x"05",x"ac"),
   841 => (x"df",x"49",x"75",x"87"),
   842 => (x"cd",x"89",x"c1",x"99"),
   843 => (x"f4",x"ec",x"c2",x"91"),
   844 => (x"4a",x"a3",x"c1",x"81"),
   845 => (x"a3",x"c3",x"51",x"12"),
   846 => (x"c5",x"51",x"12",x"4a"),
   847 => (x"51",x"12",x"4a",x"a3"),
   848 => (x"12",x"4a",x"a3",x"c7"),
   849 => (x"4a",x"a3",x"c9",x"51"),
   850 => (x"a3",x"ce",x"51",x"12"),
   851 => (x"d0",x"51",x"12",x"4a"),
   852 => (x"51",x"12",x"4a",x"a3"),
   853 => (x"12",x"4a",x"a3",x"d2"),
   854 => (x"4a",x"a3",x"d4",x"51"),
   855 => (x"a3",x"d6",x"51",x"12"),
   856 => (x"d8",x"51",x"12",x"4a"),
   857 => (x"51",x"12",x"4a",x"a3"),
   858 => (x"12",x"4a",x"a3",x"dc"),
   859 => (x"4a",x"a3",x"de",x"51"),
   860 => (x"7e",x"c1",x"51",x"12"),
   861 => (x"74",x"87",x"fc",x"c0"),
   862 => (x"05",x"99",x"c8",x"49"),
   863 => (x"74",x"87",x"ed",x"c0"),
   864 => (x"05",x"99",x"d0",x"49"),
   865 => (x"e0",x"c0",x"87",x"d3"),
   866 => (x"cc",x"c0",x"02",x"66"),
   867 => (x"c0",x"49",x"73",x"87"),
   868 => (x"70",x"0f",x"66",x"e0"),
   869 => (x"d3",x"c0",x"02",x"98"),
   870 => (x"c0",x"05",x"6e",x"87"),
   871 => (x"ec",x"c2",x"87",x"c6"),
   872 => (x"50",x"c0",x"48",x"f4"),
   873 => (x"bf",x"e8",x"f9",x"c0"),
   874 => (x"87",x"e9",x"c2",x"48"),
   875 => (x"48",x"c1",x"ed",x"c2"),
   876 => (x"c2",x"7e",x"50",x"c0"),
   877 => (x"49",x"bf",x"f0",x"ec"),
   878 => (x"bf",x"e0",x"e4",x"c2"),
   879 => (x"04",x"aa",x"71",x"4a"),
   880 => (x"cf",x"87",x"f4",x"fb"),
   881 => (x"f8",x"ff",x"ff",x"ff"),
   882 => (x"e4",x"f1",x"c2",x"4c"),
   883 => (x"c8",x"c0",x"05",x"bf"),
   884 => (x"ec",x"ec",x"c2",x"87"),
   885 => (x"fa",x"c1",x"02",x"bf"),
   886 => (x"dc",x"e4",x"c2",x"87"),
   887 => (x"c0",x"eb",x"49",x"bf"),
   888 => (x"e0",x"e4",x"c2",x"87"),
   889 => (x"48",x"a6",x"c4",x"58"),
   890 => (x"bf",x"dc",x"e4",x"c2"),
   891 => (x"ec",x"ec",x"c2",x"78"),
   892 => (x"db",x"c0",x"02",x"bf"),
   893 => (x"49",x"66",x"c4",x"87"),
   894 => (x"a9",x"74",x"99",x"74"),
   895 => (x"87",x"c8",x"c0",x"02"),
   896 => (x"c0",x"48",x"a6",x"c8"),
   897 => (x"87",x"e7",x"c0",x"78"),
   898 => (x"c1",x"48",x"a6",x"c8"),
   899 => (x"87",x"df",x"c0",x"78"),
   900 => (x"cf",x"49",x"66",x"c4"),
   901 => (x"a9",x"99",x"f8",x"ff"),
   902 => (x"87",x"c8",x"c0",x"02"),
   903 => (x"c0",x"48",x"a6",x"cc"),
   904 => (x"87",x"c5",x"c0",x"78"),
   905 => (x"c1",x"48",x"a6",x"cc"),
   906 => (x"48",x"a6",x"c8",x"78"),
   907 => (x"c8",x"78",x"66",x"cc"),
   908 => (x"de",x"c0",x"05",x"66"),
   909 => (x"49",x"66",x"c4",x"87"),
   910 => (x"ec",x"c2",x"89",x"c2"),
   911 => (x"c2",x"91",x"bf",x"e4"),
   912 => (x"48",x"bf",x"c8",x"f1"),
   913 => (x"e4",x"c2",x"80",x"71"),
   914 => (x"e4",x"c2",x"58",x"dc"),
   915 => (x"78",x"c0",x"48",x"e0"),
   916 => (x"c0",x"87",x"d4",x"f9"),
   917 => (x"ff",x"ff",x"cf",x"48"),
   918 => (x"f0",x"4c",x"f8",x"ff"),
   919 => (x"26",x"4d",x"26",x"8e"),
   920 => (x"26",x"4b",x"26",x"4c"),
   921 => (x"00",x"00",x"00",x"4f"),
   922 => (x"00",x"00",x"00",x"00"),
   923 => (x"ff",x"ff",x"ff",x"ff"),
   924 => (x"48",x"d4",x"ff",x"1e"),
   925 => (x"68",x"78",x"ff",x"c3"),
   926 => (x"1e",x"4f",x"26",x"48"),
   927 => (x"c3",x"48",x"d4",x"ff"),
   928 => (x"d0",x"ff",x"78",x"ff"),
   929 => (x"78",x"e1",x"c0",x"48"),
   930 => (x"d4",x"48",x"d4",x"ff"),
   931 => (x"1e",x"4f",x"26",x"78"),
   932 => (x"c0",x"48",x"d0",x"ff"),
   933 => (x"4f",x"26",x"78",x"e0"),
   934 => (x"87",x"d4",x"ff",x"1e"),
   935 => (x"02",x"99",x"49",x"70"),
   936 => (x"fb",x"c0",x"87",x"c6"),
   937 => (x"87",x"f1",x"05",x"a9"),
   938 => (x"4f",x"26",x"48",x"71"),
   939 => (x"5c",x"5b",x"5e",x"0e"),
   940 => (x"c0",x"4b",x"71",x"0e"),
   941 => (x"87",x"f8",x"fe",x"4c"),
   942 => (x"02",x"99",x"49",x"70"),
   943 => (x"c0",x"87",x"f9",x"c0"),
   944 => (x"c0",x"02",x"a9",x"ec"),
   945 => (x"fb",x"c0",x"87",x"f2"),
   946 => (x"eb",x"c0",x"02",x"a9"),
   947 => (x"b7",x"66",x"cc",x"87"),
   948 => (x"87",x"c7",x"03",x"ac"),
   949 => (x"c2",x"02",x"66",x"d0"),
   950 => (x"71",x"53",x"71",x"87"),
   951 => (x"87",x"c2",x"02",x"99"),
   952 => (x"cb",x"fe",x"84",x"c1"),
   953 => (x"99",x"49",x"70",x"87"),
   954 => (x"c0",x"87",x"cd",x"02"),
   955 => (x"c7",x"02",x"a9",x"ec"),
   956 => (x"a9",x"fb",x"c0",x"87"),
   957 => (x"87",x"d5",x"ff",x"05"),
   958 => (x"c3",x"02",x"66",x"d0"),
   959 => (x"7b",x"97",x"c0",x"87"),
   960 => (x"05",x"a9",x"fb",x"c0"),
   961 => (x"4a",x"74",x"87",x"c7"),
   962 => (x"c2",x"8a",x"0a",x"c0"),
   963 => (x"72",x"4a",x"74",x"87"),
   964 => (x"26",x"4c",x"26",x"48"),
   965 => (x"1e",x"4f",x"26",x"4b"),
   966 => (x"70",x"87",x"d5",x"fd"),
   967 => (x"a9",x"f0",x"c0",x"49"),
   968 => (x"c0",x"87",x"c9",x"04"),
   969 => (x"c3",x"01",x"a9",x"f9"),
   970 => (x"89",x"f0",x"c0",x"87"),
   971 => (x"04",x"a9",x"c1",x"c1"),
   972 => (x"da",x"c1",x"87",x"c9"),
   973 => (x"87",x"c3",x"01",x"a9"),
   974 => (x"71",x"89",x"f7",x"c0"),
   975 => (x"0e",x"4f",x"26",x"48"),
   976 => (x"5d",x"5c",x"5b",x"5e"),
   977 => (x"71",x"86",x"f8",x"0e"),
   978 => (x"fc",x"7e",x"c0",x"4c"),
   979 => (x"4b",x"c0",x"87",x"ed"),
   980 => (x"97",x"e0",x"ff",x"c0"),
   981 => (x"a9",x"c0",x"49",x"bf"),
   982 => (x"fc",x"87",x"cf",x"04"),
   983 => (x"83",x"c1",x"87",x"fa"),
   984 => (x"97",x"e0",x"ff",x"c0"),
   985 => (x"06",x"ab",x"49",x"bf"),
   986 => (x"ff",x"c0",x"87",x"f1"),
   987 => (x"02",x"bf",x"97",x"e0"),
   988 => (x"fb",x"fb",x"87",x"cf"),
   989 => (x"99",x"49",x"70",x"87"),
   990 => (x"c0",x"87",x"c6",x"02"),
   991 => (x"f1",x"05",x"a9",x"ec"),
   992 => (x"fb",x"4b",x"c0",x"87"),
   993 => (x"4d",x"70",x"87",x"ea"),
   994 => (x"c8",x"87",x"e5",x"fb"),
   995 => (x"df",x"fb",x"58",x"a6"),
   996 => (x"c1",x"4a",x"70",x"87"),
   997 => (x"49",x"a4",x"c8",x"83"),
   998 => (x"ad",x"49",x"69",x"97"),
   999 => (x"c9",x"87",x"da",x"05"),
  1000 => (x"69",x"97",x"49",x"a4"),
  1001 => (x"a9",x"66",x"c4",x"49"),
  1002 => (x"ca",x"87",x"ce",x"05"),
  1003 => (x"69",x"97",x"49",x"a4"),
  1004 => (x"c4",x"05",x"aa",x"49"),
  1005 => (x"d0",x"7e",x"c1",x"87"),
  1006 => (x"ad",x"ec",x"c0",x"87"),
  1007 => (x"c0",x"87",x"c6",x"02"),
  1008 => (x"c4",x"05",x"ad",x"fb"),
  1009 => (x"c1",x"4b",x"c0",x"87"),
  1010 => (x"fe",x"02",x"6e",x"7e"),
  1011 => (x"fe",x"fa",x"87",x"f5"),
  1012 => (x"f8",x"48",x"73",x"87"),
  1013 => (x"26",x"4d",x"26",x"8e"),
  1014 => (x"26",x"4b",x"26",x"4c"),
  1015 => (x"00",x"00",x"00",x"4f"),
  1016 => (x"1e",x"73",x"1e",x"00"),
  1017 => (x"c8",x"4b",x"d4",x"ff"),
  1018 => (x"d0",x"ff",x"4a",x"66"),
  1019 => (x"78",x"c5",x"c8",x"48"),
  1020 => (x"c1",x"48",x"d4",x"ff"),
  1021 => (x"7b",x"11",x"78",x"d4"),
  1022 => (x"f9",x"05",x"8a",x"c1"),
  1023 => (x"48",x"d0",x"ff",x"87"),
  1024 => (x"4b",x"26",x"78",x"c4"),
  1025 => (x"5e",x"0e",x"4f",x"26"),
  1026 => (x"0e",x"5d",x"5c",x"5b"),
  1027 => (x"7e",x"71",x"86",x"f8"),
  1028 => (x"f1",x"c2",x"1e",x"6e"),
  1029 => (x"ff",x"e3",x"49",x"f8"),
  1030 => (x"70",x"86",x"c4",x"87"),
  1031 => (x"e4",x"c4",x"02",x"98"),
  1032 => (x"c8",x"ed",x"c1",x"87"),
  1033 => (x"49",x"6e",x"4c",x"bf"),
  1034 => (x"c8",x"87",x"d4",x"fc"),
  1035 => (x"98",x"70",x"58",x"a6"),
  1036 => (x"c4",x"87",x"c5",x"05"),
  1037 => (x"78",x"c1",x"48",x"a6"),
  1038 => (x"c5",x"48",x"d0",x"ff"),
  1039 => (x"48",x"d4",x"ff",x"78"),
  1040 => (x"c4",x"78",x"d5",x"c1"),
  1041 => (x"89",x"c1",x"49",x"66"),
  1042 => (x"ed",x"c1",x"31",x"c6"),
  1043 => (x"4a",x"bf",x"97",x"c0"),
  1044 => (x"ff",x"b0",x"71",x"48"),
  1045 => (x"ff",x"78",x"08",x"d4"),
  1046 => (x"78",x"c4",x"48",x"d0"),
  1047 => (x"97",x"f4",x"f1",x"c2"),
  1048 => (x"99",x"d0",x"49",x"bf"),
  1049 => (x"c5",x"87",x"dd",x"02"),
  1050 => (x"48",x"d4",x"ff",x"78"),
  1051 => (x"c0",x"78",x"d6",x"c1"),
  1052 => (x"48",x"d4",x"ff",x"4a"),
  1053 => (x"c1",x"78",x"ff",x"c3"),
  1054 => (x"aa",x"e0",x"c0",x"82"),
  1055 => (x"ff",x"87",x"f2",x"04"),
  1056 => (x"78",x"c4",x"48",x"d0"),
  1057 => (x"c3",x"48",x"d4",x"ff"),
  1058 => (x"d0",x"ff",x"78",x"ff"),
  1059 => (x"ff",x"78",x"c5",x"48"),
  1060 => (x"d3",x"c1",x"48",x"d4"),
  1061 => (x"ff",x"78",x"c1",x"78"),
  1062 => (x"78",x"c4",x"48",x"d0"),
  1063 => (x"06",x"ac",x"b7",x"c0"),
  1064 => (x"c2",x"87",x"cb",x"c2"),
  1065 => (x"4b",x"bf",x"c0",x"f2"),
  1066 => (x"73",x"7e",x"74",x"8c"),
  1067 => (x"dd",x"c1",x"02",x"9b"),
  1068 => (x"4d",x"c0",x"c8",x"87"),
  1069 => (x"ab",x"b7",x"c0",x"8b"),
  1070 => (x"c8",x"87",x"c6",x"03"),
  1071 => (x"c0",x"4d",x"a3",x"c0"),
  1072 => (x"f4",x"f1",x"c2",x"4b"),
  1073 => (x"d0",x"49",x"bf",x"97"),
  1074 => (x"87",x"cf",x"02",x"99"),
  1075 => (x"f1",x"c2",x"1e",x"c0"),
  1076 => (x"f7",x"e5",x"49",x"f8"),
  1077 => (x"70",x"86",x"c4",x"87"),
  1078 => (x"c2",x"87",x"d8",x"4c"),
  1079 => (x"c2",x"1e",x"e4",x"e4"),
  1080 => (x"e5",x"49",x"f8",x"f1"),
  1081 => (x"4c",x"70",x"87",x"e6"),
  1082 => (x"e4",x"c2",x"1e",x"75"),
  1083 => (x"f0",x"fb",x"49",x"e4"),
  1084 => (x"74",x"86",x"c8",x"87"),
  1085 => (x"87",x"c5",x"05",x"9c"),
  1086 => (x"ca",x"c1",x"48",x"c0"),
  1087 => (x"c2",x"1e",x"c1",x"87"),
  1088 => (x"e3",x"49",x"f8",x"f1"),
  1089 => (x"86",x"c4",x"87",x"f9"),
  1090 => (x"fe",x"05",x"9b",x"73"),
  1091 => (x"4c",x"6e",x"87",x"e3"),
  1092 => (x"06",x"ac",x"b7",x"c0"),
  1093 => (x"f1",x"c2",x"87",x"d1"),
  1094 => (x"78",x"c0",x"48",x"f8"),
  1095 => (x"78",x"c0",x"80",x"d0"),
  1096 => (x"f2",x"c2",x"80",x"f4"),
  1097 => (x"c0",x"78",x"bf",x"c4"),
  1098 => (x"fd",x"01",x"ac",x"b7"),
  1099 => (x"d0",x"ff",x"87",x"f5"),
  1100 => (x"ff",x"78",x"c5",x"48"),
  1101 => (x"d3",x"c1",x"48",x"d4"),
  1102 => (x"ff",x"78",x"c0",x"78"),
  1103 => (x"78",x"c4",x"48",x"d0"),
  1104 => (x"c2",x"c0",x"48",x"c1"),
  1105 => (x"f8",x"48",x"c0",x"87"),
  1106 => (x"26",x"4d",x"26",x"8e"),
  1107 => (x"26",x"4b",x"26",x"4c"),
  1108 => (x"5b",x"5e",x"0e",x"4f"),
  1109 => (x"fc",x"0e",x"5d",x"5c"),
  1110 => (x"c0",x"4d",x"71",x"86"),
  1111 => (x"04",x"ad",x"4c",x"4b"),
  1112 => (x"c0",x"87",x"e8",x"c0"),
  1113 => (x"74",x"1e",x"ff",x"fc"),
  1114 => (x"87",x"c4",x"02",x"9c"),
  1115 => (x"87",x"c2",x"4a",x"c0"),
  1116 => (x"49",x"72",x"4a",x"c1"),
  1117 => (x"c4",x"87",x"fa",x"eb"),
  1118 => (x"c1",x"7e",x"70",x"86"),
  1119 => (x"c2",x"05",x"6e",x"83"),
  1120 => (x"c1",x"4b",x"75",x"87"),
  1121 => (x"06",x"ab",x"75",x"84"),
  1122 => (x"6e",x"87",x"d8",x"ff"),
  1123 => (x"26",x"8e",x"fc",x"48"),
  1124 => (x"26",x"4c",x"26",x"4d"),
  1125 => (x"0e",x"4f",x"26",x"4b"),
  1126 => (x"0e",x"5c",x"5b",x"5e"),
  1127 => (x"66",x"cc",x"4b",x"71"),
  1128 => (x"4c",x"87",x"d8",x"02"),
  1129 => (x"02",x"8c",x"f0",x"c0"),
  1130 => (x"4a",x"74",x"87",x"d8"),
  1131 => (x"d1",x"02",x"8a",x"c1"),
  1132 => (x"cd",x"02",x"8a",x"87"),
  1133 => (x"c9",x"02",x"8a",x"87"),
  1134 => (x"73",x"87",x"d9",x"87"),
  1135 => (x"87",x"c6",x"f9",x"49"),
  1136 => (x"1e",x"74",x"87",x"d2"),
  1137 => (x"d9",x"c1",x"49",x"c0"),
  1138 => (x"1e",x"74",x"87",x"de"),
  1139 => (x"d9",x"c1",x"49",x"73"),
  1140 => (x"86",x"c8",x"87",x"d6"),
  1141 => (x"4b",x"26",x"4c",x"26"),
  1142 => (x"5e",x"0e",x"4f",x"26"),
  1143 => (x"0e",x"5d",x"5c",x"5b"),
  1144 => (x"4c",x"71",x"86",x"fc"),
  1145 => (x"c2",x"91",x"de",x"49"),
  1146 => (x"71",x"4d",x"d8",x"f3"),
  1147 => (x"02",x"6d",x"97",x"85"),
  1148 => (x"c2",x"87",x"dc",x"c1"),
  1149 => (x"49",x"bf",x"c8",x"f3"),
  1150 => (x"fd",x"71",x"81",x"74"),
  1151 => (x"7e",x"70",x"87",x"d3"),
  1152 => (x"c0",x"02",x"98",x"48"),
  1153 => (x"f3",x"c2",x"87",x"f2"),
  1154 => (x"4a",x"70",x"4b",x"cc"),
  1155 => (x"fb",x"fe",x"49",x"cb"),
  1156 => (x"4b",x"74",x"87",x"ee"),
  1157 => (x"ed",x"c1",x"93",x"cc"),
  1158 => (x"83",x"c4",x"83",x"cc"),
  1159 => (x"7b",x"dc",x"c9",x"c1"),
  1160 => (x"c2",x"c1",x"49",x"74"),
  1161 => (x"7b",x"75",x"87",x"fa"),
  1162 => (x"97",x"c4",x"ed",x"c1"),
  1163 => (x"c2",x"1e",x"49",x"bf"),
  1164 => (x"fd",x"49",x"cc",x"f3"),
  1165 => (x"86",x"c4",x"87",x"e1"),
  1166 => (x"c2",x"c1",x"49",x"74"),
  1167 => (x"49",x"c0",x"87",x"e2"),
  1168 => (x"87",x"fd",x"c3",x"c1"),
  1169 => (x"48",x"f0",x"f1",x"c2"),
  1170 => (x"c0",x"49",x"50",x"c0"),
  1171 => (x"fc",x"87",x"c3",x"e1"),
  1172 => (x"26",x"4d",x"26",x"8e"),
  1173 => (x"26",x"4b",x"26",x"4c"),
  1174 => (x"00",x"00",x"00",x"4f"),
  1175 => (x"64",x"61",x"6f",x"4c"),
  1176 => (x"2e",x"67",x"6e",x"69"),
  1177 => (x"00",x"00",x"2e",x"2e"),
  1178 => (x"61",x"42",x"20",x"80"),
  1179 => (x"00",x"00",x"6b",x"63"),
  1180 => (x"64",x"61",x"6f",x"4c"),
  1181 => (x"20",x"2e",x"2a",x"20"),
  1182 => (x"00",x"00",x"00",x"00"),
  1183 => (x"00",x"00",x"20",x"3a"),
  1184 => (x"61",x"42",x"20",x"80"),
  1185 => (x"00",x"00",x"6b",x"63"),
  1186 => (x"78",x"45",x"20",x"80"),
  1187 => (x"00",x"00",x"74",x"69"),
  1188 => (x"49",x"20",x"44",x"53"),
  1189 => (x"2e",x"74",x"69",x"6e"),
  1190 => (x"00",x"00",x"00",x"2e"),
  1191 => (x"00",x"00",x"4b",x"4f"),
  1192 => (x"54",x"4f",x"4f",x"42"),
  1193 => (x"20",x"20",x"20",x"20"),
  1194 => (x"00",x"4d",x"4f",x"52"),
  1195 => (x"71",x"1e",x"73",x"1e"),
  1196 => (x"f3",x"c2",x"49",x"4b"),
  1197 => (x"71",x"81",x"bf",x"c8"),
  1198 => (x"70",x"87",x"d6",x"fa"),
  1199 => (x"c4",x"02",x"9a",x"4a"),
  1200 => (x"e6",x"e4",x"49",x"87"),
  1201 => (x"c8",x"f3",x"c2",x"87"),
  1202 => (x"73",x"78",x"c0",x"48"),
  1203 => (x"87",x"fa",x"c1",x"49"),
  1204 => (x"4f",x"26",x"4b",x"26"),
  1205 => (x"71",x"1e",x"73",x"1e"),
  1206 => (x"4a",x"a3",x"c4",x"4b"),
  1207 => (x"87",x"d0",x"c1",x"02"),
  1208 => (x"dc",x"02",x"8a",x"c1"),
  1209 => (x"c0",x"02",x"8a",x"87"),
  1210 => (x"05",x"8a",x"87",x"f2"),
  1211 => (x"c2",x"87",x"d3",x"c1"),
  1212 => (x"02",x"bf",x"c8",x"f3"),
  1213 => (x"48",x"87",x"cb",x"c1"),
  1214 => (x"f3",x"c2",x"88",x"c1"),
  1215 => (x"c1",x"c1",x"58",x"cc"),
  1216 => (x"c8",x"f3",x"c2",x"87"),
  1217 => (x"89",x"c6",x"49",x"bf"),
  1218 => (x"59",x"cc",x"f3",x"c2"),
  1219 => (x"03",x"a9",x"b7",x"c0"),
  1220 => (x"c2",x"87",x"ef",x"c0"),
  1221 => (x"c0",x"48",x"c8",x"f3"),
  1222 => (x"87",x"e6",x"c0",x"78"),
  1223 => (x"bf",x"c4",x"f3",x"c2"),
  1224 => (x"c2",x"87",x"df",x"02"),
  1225 => (x"48",x"bf",x"c8",x"f3"),
  1226 => (x"f3",x"c2",x"80",x"c1"),
  1227 => (x"87",x"d2",x"58",x"cc"),
  1228 => (x"bf",x"c4",x"f3",x"c2"),
  1229 => (x"c2",x"87",x"cb",x"02"),
  1230 => (x"48",x"bf",x"c8",x"f3"),
  1231 => (x"f3",x"c2",x"80",x"c6"),
  1232 => (x"49",x"73",x"58",x"cc"),
  1233 => (x"4b",x"26",x"87",x"c4"),
  1234 => (x"5e",x"0e",x"4f",x"26"),
  1235 => (x"0e",x"5d",x"5c",x"5b"),
  1236 => (x"a6",x"d0",x"86",x"f0"),
  1237 => (x"e4",x"e4",x"c2",x"59"),
  1238 => (x"c2",x"4c",x"c0",x"4d"),
  1239 => (x"c1",x"48",x"c4",x"f3"),
  1240 => (x"48",x"a6",x"c8",x"78"),
  1241 => (x"7e",x"75",x"78",x"c0"),
  1242 => (x"bf",x"c8",x"f3",x"c2"),
  1243 => (x"06",x"a8",x"c0",x"48"),
  1244 => (x"c8",x"87",x"c0",x"c1"),
  1245 => (x"7e",x"75",x"5c",x"a6"),
  1246 => (x"48",x"e4",x"e4",x"c2"),
  1247 => (x"f2",x"c0",x"02",x"98"),
  1248 => (x"4d",x"66",x"c4",x"87"),
  1249 => (x"1e",x"ff",x"fc",x"c0"),
  1250 => (x"c4",x"02",x"66",x"cc"),
  1251 => (x"c2",x"4c",x"c0",x"87"),
  1252 => (x"74",x"4c",x"c1",x"87"),
  1253 => (x"87",x"d9",x"e3",x"49"),
  1254 => (x"7e",x"70",x"86",x"c4"),
  1255 => (x"66",x"c8",x"85",x"c1"),
  1256 => (x"cc",x"80",x"c1",x"48"),
  1257 => (x"f3",x"c2",x"58",x"a6"),
  1258 => (x"03",x"ad",x"bf",x"c8"),
  1259 => (x"05",x"6e",x"87",x"c5"),
  1260 => (x"6e",x"87",x"d1",x"ff"),
  1261 => (x"75",x"4c",x"c0",x"4d"),
  1262 => (x"dc",x"c3",x"02",x"9d"),
  1263 => (x"ff",x"fc",x"c0",x"87"),
  1264 => (x"02",x"66",x"cc",x"1e"),
  1265 => (x"a6",x"c8",x"87",x"c7"),
  1266 => (x"c5",x"78",x"c0",x"48"),
  1267 => (x"48",x"a6",x"c8",x"87"),
  1268 => (x"66",x"c8",x"78",x"c1"),
  1269 => (x"87",x"d9",x"e2",x"49"),
  1270 => (x"7e",x"70",x"86",x"c4"),
  1271 => (x"c2",x"02",x"98",x"48"),
  1272 => (x"cb",x"49",x"87",x"e4"),
  1273 => (x"49",x"69",x"97",x"81"),
  1274 => (x"c1",x"02",x"99",x"d0"),
  1275 => (x"49",x"74",x"87",x"d4"),
  1276 => (x"ed",x"c1",x"91",x"cc"),
  1277 => (x"ca",x"c1",x"81",x"cc"),
  1278 => (x"81",x"c8",x"79",x"ec"),
  1279 => (x"74",x"51",x"ff",x"c3"),
  1280 => (x"c2",x"91",x"de",x"49"),
  1281 => (x"71",x"4d",x"d8",x"f3"),
  1282 => (x"97",x"c1",x"c2",x"85"),
  1283 => (x"49",x"a5",x"c1",x"7d"),
  1284 => (x"c2",x"51",x"e0",x"c0"),
  1285 => (x"bf",x"97",x"f4",x"ec"),
  1286 => (x"c1",x"87",x"d2",x"02"),
  1287 => (x"4b",x"a5",x"c2",x"84"),
  1288 => (x"4a",x"f4",x"ec",x"c2"),
  1289 => (x"f3",x"fe",x"49",x"db"),
  1290 => (x"d9",x"c1",x"87",x"d6"),
  1291 => (x"49",x"a5",x"cd",x"87"),
  1292 => (x"84",x"c1",x"51",x"c0"),
  1293 => (x"6e",x"4b",x"a5",x"c2"),
  1294 => (x"fe",x"49",x"cb",x"4a"),
  1295 => (x"c1",x"87",x"c1",x"f3"),
  1296 => (x"49",x"74",x"87",x"c4"),
  1297 => (x"ed",x"c1",x"91",x"cc"),
  1298 => (x"c7",x"c1",x"81",x"cc"),
  1299 => (x"ec",x"c2",x"79",x"da"),
  1300 => (x"02",x"bf",x"97",x"f4"),
  1301 => (x"49",x"74",x"87",x"d8"),
  1302 => (x"84",x"c1",x"91",x"de"),
  1303 => (x"4b",x"d8",x"f3",x"c2"),
  1304 => (x"ec",x"c2",x"83",x"71"),
  1305 => (x"49",x"dd",x"4a",x"f4"),
  1306 => (x"87",x"d4",x"f2",x"fe"),
  1307 => (x"4b",x"74",x"87",x"d8"),
  1308 => (x"f3",x"c2",x"93",x"de"),
  1309 => (x"a3",x"cb",x"83",x"d8"),
  1310 => (x"c1",x"51",x"c0",x"49"),
  1311 => (x"4a",x"6e",x"73",x"84"),
  1312 => (x"f1",x"fe",x"49",x"cb"),
  1313 => (x"66",x"c8",x"87",x"fa"),
  1314 => (x"cc",x"80",x"c1",x"48"),
  1315 => (x"ac",x"c7",x"58",x"a6"),
  1316 => (x"87",x"c5",x"c0",x"03"),
  1317 => (x"e4",x"fc",x"05",x"6e"),
  1318 => (x"03",x"ac",x"c7",x"87"),
  1319 => (x"c2",x"87",x"e4",x"c0"),
  1320 => (x"c0",x"48",x"c4",x"f3"),
  1321 => (x"cc",x"49",x"74",x"78"),
  1322 => (x"cc",x"ed",x"c1",x"91"),
  1323 => (x"da",x"c7",x"c1",x"81"),
  1324 => (x"de",x"49",x"74",x"79"),
  1325 => (x"d8",x"f3",x"c2",x"91"),
  1326 => (x"c1",x"51",x"c0",x"81"),
  1327 => (x"04",x"ac",x"c7",x"84"),
  1328 => (x"c1",x"87",x"dc",x"ff"),
  1329 => (x"c0",x"48",x"e8",x"ee"),
  1330 => (x"c1",x"80",x"f7",x"50"),
  1331 => (x"c1",x"40",x"f0",x"d4"),
  1332 => (x"c8",x"78",x"e8",x"c9"),
  1333 => (x"d4",x"cb",x"c1",x"80"),
  1334 => (x"49",x"66",x"cc",x"78"),
  1335 => (x"87",x"c0",x"f8",x"c0"),
  1336 => (x"4d",x"26",x"8e",x"f0"),
  1337 => (x"4b",x"26",x"4c",x"26"),
  1338 => (x"73",x"1e",x"4f",x"26"),
  1339 => (x"49",x"4b",x"71",x"1e"),
  1340 => (x"ed",x"c1",x"91",x"cc"),
  1341 => (x"a1",x"c8",x"81",x"cc"),
  1342 => (x"c0",x"ed",x"c1",x"4a"),
  1343 => (x"c9",x"50",x"12",x"48"),
  1344 => (x"ff",x"c0",x"4a",x"a1"),
  1345 => (x"50",x"12",x"48",x"e0"),
  1346 => (x"ed",x"c1",x"81",x"ca"),
  1347 => (x"50",x"11",x"48",x"c4"),
  1348 => (x"97",x"c4",x"ed",x"c1"),
  1349 => (x"c0",x"1e",x"49",x"bf"),
  1350 => (x"87",x"fb",x"f1",x"49"),
  1351 => (x"e9",x"f8",x"49",x"73"),
  1352 => (x"26",x"8e",x"fc",x"87"),
  1353 => (x"1e",x"4f",x"26",x"4b"),
  1354 => (x"f8",x"c0",x"49",x"c0"),
  1355 => (x"4f",x"26",x"87",x"d3"),
  1356 => (x"49",x"4a",x"71",x"1e"),
  1357 => (x"ed",x"c1",x"91",x"cc"),
  1358 => (x"81",x"c8",x"81",x"cc"),
  1359 => (x"48",x"f0",x"f1",x"c2"),
  1360 => (x"f0",x"c0",x"50",x"11"),
  1361 => (x"ed",x"fe",x"49",x"a2"),
  1362 => (x"49",x"c0",x"87",x"c2"),
  1363 => (x"26",x"87",x"c3",x"d5"),
  1364 => (x"d4",x"ff",x"1e",x"4f"),
  1365 => (x"7a",x"ff",x"c3",x"4a"),
  1366 => (x"c0",x"48",x"d0",x"ff"),
  1367 => (x"7a",x"de",x"78",x"e1"),
  1368 => (x"c8",x"48",x"7a",x"71"),
  1369 => (x"7a",x"70",x"28",x"b7"),
  1370 => (x"b7",x"d0",x"48",x"71"),
  1371 => (x"71",x"7a",x"70",x"28"),
  1372 => (x"28",x"b7",x"d8",x"48"),
  1373 => (x"d0",x"ff",x"7a",x"70"),
  1374 => (x"78",x"e0",x"c0",x"48"),
  1375 => (x"5e",x"0e",x"4f",x"26"),
  1376 => (x"0e",x"5d",x"5c",x"5b"),
  1377 => (x"4d",x"71",x"86",x"f4"),
  1378 => (x"c1",x"91",x"cc",x"49"),
  1379 => (x"c8",x"81",x"cc",x"ed"),
  1380 => (x"a1",x"ca",x"4a",x"a1"),
  1381 => (x"48",x"a6",x"c4",x"7e"),
  1382 => (x"bf",x"ec",x"f1",x"c2"),
  1383 => (x"bf",x"97",x"6e",x"78"),
  1384 => (x"4c",x"66",x"c4",x"4b"),
  1385 => (x"48",x"12",x"2c",x"73"),
  1386 => (x"70",x"58",x"a6",x"cc"),
  1387 => (x"c9",x"84",x"c1",x"9c"),
  1388 => (x"49",x"69",x"97",x"81"),
  1389 => (x"c2",x"04",x"ac",x"b7"),
  1390 => (x"6e",x"4c",x"c0",x"87"),
  1391 => (x"c8",x"4a",x"bf",x"97"),
  1392 => (x"31",x"72",x"49",x"66"),
  1393 => (x"66",x"c4",x"b9",x"ff"),
  1394 => (x"72",x"48",x"74",x"99"),
  1395 => (x"b1",x"4a",x"70",x"30"),
  1396 => (x"59",x"f0",x"f1",x"c2"),
  1397 => (x"87",x"f9",x"fd",x"71"),
  1398 => (x"f3",x"c2",x"1e",x"c7"),
  1399 => (x"c1",x"1e",x"bf",x"c0"),
  1400 => (x"c2",x"1e",x"cc",x"ed"),
  1401 => (x"bf",x"97",x"f0",x"f1"),
  1402 => (x"87",x"f4",x"c1",x"49"),
  1403 => (x"f3",x"c0",x"49",x"75"),
  1404 => (x"8e",x"e8",x"87",x"ee"),
  1405 => (x"4c",x"26",x"4d",x"26"),
  1406 => (x"4f",x"26",x"4b",x"26"),
  1407 => (x"71",x"1e",x"73",x"1e"),
  1408 => (x"f9",x"fd",x"49",x"4b"),
  1409 => (x"fd",x"49",x"73",x"87"),
  1410 => (x"4b",x"26",x"87",x"f4"),
  1411 => (x"73",x"1e",x"4f",x"26"),
  1412 => (x"c2",x"4b",x"71",x"1e"),
  1413 => (x"d6",x"02",x"4a",x"a3"),
  1414 => (x"05",x"8a",x"c1",x"87"),
  1415 => (x"c2",x"87",x"e2",x"c0"),
  1416 => (x"02",x"bf",x"c0",x"f3"),
  1417 => (x"c1",x"48",x"87",x"db"),
  1418 => (x"c4",x"f3",x"c2",x"88"),
  1419 => (x"c2",x"87",x"d2",x"58"),
  1420 => (x"02",x"bf",x"c4",x"f3"),
  1421 => (x"f3",x"c2",x"87",x"cb"),
  1422 => (x"c1",x"48",x"bf",x"c0"),
  1423 => (x"c4",x"f3",x"c2",x"80"),
  1424 => (x"c2",x"1e",x"c7",x"58"),
  1425 => (x"1e",x"bf",x"c0",x"f3"),
  1426 => (x"1e",x"cc",x"ed",x"c1"),
  1427 => (x"97",x"f0",x"f1",x"c2"),
  1428 => (x"87",x"cc",x"49",x"bf"),
  1429 => (x"f2",x"c0",x"49",x"73"),
  1430 => (x"8e",x"f4",x"87",x"c6"),
  1431 => (x"4f",x"26",x"4b",x"26"),
  1432 => (x"5c",x"5b",x"5e",x"0e"),
  1433 => (x"cc",x"ff",x"0e",x"5d"),
  1434 => (x"a6",x"e8",x"c0",x"86"),
  1435 => (x"48",x"a6",x"cc",x"59"),
  1436 => (x"80",x"c4",x"78",x"c0"),
  1437 => (x"80",x"c4",x"78",x"c0"),
  1438 => (x"80",x"c4",x"78",x"c0"),
  1439 => (x"78",x"66",x"c8",x"c1"),
  1440 => (x"78",x"c1",x"80",x"c4"),
  1441 => (x"78",x"c1",x"80",x"c4"),
  1442 => (x"48",x"c4",x"f3",x"c2"),
  1443 => (x"df",x"ff",x"78",x"c1"),
  1444 => (x"c3",x"e0",x"87",x"e9"),
  1445 => (x"d7",x"df",x"ff",x"87"),
  1446 => (x"c0",x"4d",x"70",x"87"),
  1447 => (x"c1",x"02",x"ad",x"fb"),
  1448 => (x"e4",x"c0",x"87",x"f3"),
  1449 => (x"e8",x"c1",x"05",x"66"),
  1450 => (x"66",x"c4",x"c1",x"87"),
  1451 => (x"6a",x"82",x"c4",x"4a"),
  1452 => (x"f0",x"c9",x"c1",x"7e"),
  1453 => (x"20",x"49",x"6e",x"48"),
  1454 => (x"10",x"41",x"20",x"41"),
  1455 => (x"66",x"c4",x"c1",x"51"),
  1456 => (x"ea",x"d3",x"c1",x"48"),
  1457 => (x"c7",x"49",x"6a",x"78"),
  1458 => (x"c1",x"51",x"75",x"81"),
  1459 => (x"c8",x"49",x"66",x"c4"),
  1460 => (x"dc",x"51",x"c1",x"81"),
  1461 => (x"78",x"c2",x"48",x"a6"),
  1462 => (x"49",x"66",x"c4",x"c1"),
  1463 => (x"51",x"c0",x"81",x"c9"),
  1464 => (x"49",x"66",x"c4",x"c1"),
  1465 => (x"51",x"c0",x"81",x"ca"),
  1466 => (x"1e",x"d8",x"1e",x"c1"),
  1467 => (x"81",x"c8",x"49",x"6a"),
  1468 => (x"87",x"f8",x"de",x"ff"),
  1469 => (x"c8",x"c1",x"86",x"c8"),
  1470 => (x"a8",x"c0",x"48",x"66"),
  1471 => (x"d4",x"87",x"c7",x"01"),
  1472 => (x"78",x"c1",x"48",x"a6"),
  1473 => (x"c8",x"c1",x"87",x"cf"),
  1474 => (x"88",x"c1",x"48",x"66"),
  1475 => (x"c4",x"58",x"a6",x"dc"),
  1476 => (x"c3",x"de",x"ff",x"87"),
  1477 => (x"02",x"9d",x"75",x"87"),
  1478 => (x"d4",x"87",x"f1",x"cb"),
  1479 => (x"cc",x"c1",x"48",x"66"),
  1480 => (x"cb",x"03",x"a8",x"66"),
  1481 => (x"7e",x"c0",x"87",x"e6"),
  1482 => (x"87",x"c4",x"dd",x"ff"),
  1483 => (x"c1",x"48",x"4d",x"70"),
  1484 => (x"a6",x"c8",x"88",x"c6"),
  1485 => (x"02",x"98",x"70",x"58"),
  1486 => (x"48",x"87",x"d6",x"c1"),
  1487 => (x"a6",x"c8",x"88",x"c9"),
  1488 => (x"02",x"98",x"70",x"58"),
  1489 => (x"48",x"87",x"d7",x"c5"),
  1490 => (x"a6",x"c8",x"88",x"c1"),
  1491 => (x"02",x"98",x"70",x"58"),
  1492 => (x"48",x"87",x"f8",x"c2"),
  1493 => (x"a6",x"c8",x"88",x"c3"),
  1494 => (x"02",x"98",x"70",x"58"),
  1495 => (x"c1",x"48",x"87",x"cf"),
  1496 => (x"58",x"a6",x"c8",x"88"),
  1497 => (x"c4",x"02",x"98",x"70"),
  1498 => (x"fe",x"c9",x"87",x"f4"),
  1499 => (x"7e",x"f0",x"c0",x"87"),
  1500 => (x"87",x"fc",x"db",x"ff"),
  1501 => (x"ec",x"c0",x"4d",x"70"),
  1502 => (x"87",x"c2",x"02",x"ad"),
  1503 => (x"ec",x"c0",x"7e",x"75"),
  1504 => (x"87",x"cd",x"02",x"ad"),
  1505 => (x"87",x"e8",x"db",x"ff"),
  1506 => (x"ec",x"c0",x"4d",x"70"),
  1507 => (x"f3",x"ff",x"05",x"ad"),
  1508 => (x"66",x"e4",x"c0",x"87"),
  1509 => (x"87",x"ea",x"c1",x"05"),
  1510 => (x"02",x"ad",x"ec",x"c0"),
  1511 => (x"db",x"ff",x"87",x"c4"),
  1512 => (x"1e",x"c0",x"87",x"ce"),
  1513 => (x"66",x"dc",x"1e",x"ca"),
  1514 => (x"c1",x"93",x"cc",x"4b"),
  1515 => (x"c4",x"83",x"66",x"cc"),
  1516 => (x"49",x"6c",x"4c",x"a3"),
  1517 => (x"87",x"f4",x"db",x"ff"),
  1518 => (x"1e",x"de",x"1e",x"c1"),
  1519 => (x"db",x"ff",x"49",x"6c"),
  1520 => (x"86",x"d0",x"87",x"ea"),
  1521 => (x"7b",x"ea",x"d3",x"c1"),
  1522 => (x"dc",x"49",x"a3",x"c8"),
  1523 => (x"a3",x"c9",x"51",x"66"),
  1524 => (x"66",x"e0",x"c0",x"49"),
  1525 => (x"49",x"a3",x"ca",x"51"),
  1526 => (x"66",x"dc",x"51",x"6e"),
  1527 => (x"c0",x"80",x"c1",x"48"),
  1528 => (x"d4",x"58",x"a6",x"e0"),
  1529 => (x"66",x"d8",x"48",x"66"),
  1530 => (x"87",x"cb",x"04",x"a8"),
  1531 => (x"c1",x"48",x"66",x"d4"),
  1532 => (x"58",x"a6",x"d8",x"80"),
  1533 => (x"d8",x"87",x"fa",x"c7"),
  1534 => (x"88",x"c1",x"48",x"66"),
  1535 => (x"c7",x"58",x"a6",x"dc"),
  1536 => (x"da",x"ff",x"87",x"ef"),
  1537 => (x"4d",x"70",x"87",x"d2"),
  1538 => (x"ff",x"87",x"e6",x"c7"),
  1539 => (x"d0",x"87",x"c8",x"dc"),
  1540 => (x"66",x"d0",x"58",x"a6"),
  1541 => (x"87",x"c6",x"06",x"a8"),
  1542 => (x"cc",x"48",x"a6",x"d0"),
  1543 => (x"db",x"ff",x"78",x"66"),
  1544 => (x"ec",x"c0",x"87",x"f5"),
  1545 => (x"f5",x"c1",x"05",x"a8"),
  1546 => (x"66",x"e4",x"c0",x"87"),
  1547 => (x"87",x"e5",x"c1",x"05"),
  1548 => (x"cc",x"49",x"66",x"d4"),
  1549 => (x"66",x"c4",x"c1",x"91"),
  1550 => (x"4a",x"a1",x"c4",x"81"),
  1551 => (x"a1",x"c8",x"4c",x"6a"),
  1552 => (x"52",x"66",x"cc",x"4a"),
  1553 => (x"79",x"f0",x"d4",x"c1"),
  1554 => (x"87",x"e4",x"d8",x"ff"),
  1555 => (x"02",x"9d",x"4d",x"70"),
  1556 => (x"fb",x"c0",x"87",x"da"),
  1557 => (x"87",x"d4",x"02",x"ad"),
  1558 => (x"d8",x"ff",x"54",x"75"),
  1559 => (x"4d",x"70",x"87",x"d2"),
  1560 => (x"c7",x"c0",x"02",x"9d"),
  1561 => (x"ad",x"fb",x"c0",x"87"),
  1562 => (x"87",x"ec",x"ff",x"05"),
  1563 => (x"c2",x"54",x"e0",x"c0"),
  1564 => (x"97",x"c0",x"54",x"c1"),
  1565 => (x"48",x"66",x"d4",x"7c"),
  1566 => (x"04",x"a8",x"66",x"d8"),
  1567 => (x"d4",x"87",x"cb",x"c0"),
  1568 => (x"80",x"c1",x"48",x"66"),
  1569 => (x"c5",x"58",x"a6",x"d8"),
  1570 => (x"66",x"d8",x"87",x"e7"),
  1571 => (x"dc",x"88",x"c1",x"48"),
  1572 => (x"dc",x"c5",x"58",x"a6"),
  1573 => (x"ff",x"d7",x"ff",x"87"),
  1574 => (x"c5",x"4d",x"70",x"87"),
  1575 => (x"66",x"cc",x"87",x"d3"),
  1576 => (x"66",x"e4",x"c0",x"48"),
  1577 => (x"f4",x"c4",x"05",x"a8"),
  1578 => (x"a6",x"e8",x"c0",x"87"),
  1579 => (x"ff",x"78",x"c0",x"48"),
  1580 => (x"70",x"87",x"e4",x"d9"),
  1581 => (x"de",x"d9",x"ff",x"7e"),
  1582 => (x"a6",x"f0",x"c0",x"87"),
  1583 => (x"a8",x"ec",x"c0",x"58"),
  1584 => (x"87",x"c7",x"c0",x"05"),
  1585 => (x"78",x"6e",x"48",x"a6"),
  1586 => (x"ff",x"87",x"c4",x"c0"),
  1587 => (x"d4",x"87",x"e1",x"d6"),
  1588 => (x"91",x"cc",x"49",x"66"),
  1589 => (x"48",x"66",x"c4",x"c1"),
  1590 => (x"a6",x"c8",x"80",x"71"),
  1591 => (x"4a",x"66",x"c4",x"58"),
  1592 => (x"66",x"c4",x"82",x"c8"),
  1593 => (x"6e",x"81",x"ca",x"49"),
  1594 => (x"66",x"ec",x"c0",x"51"),
  1595 => (x"6e",x"81",x"c1",x"49"),
  1596 => (x"71",x"48",x"c1",x"89"),
  1597 => (x"c1",x"49",x"70",x"30"),
  1598 => (x"7a",x"97",x"71",x"89"),
  1599 => (x"bf",x"ec",x"f1",x"c2"),
  1600 => (x"97",x"29",x"6e",x"49"),
  1601 => (x"71",x"48",x"4a",x"6a"),
  1602 => (x"a6",x"f4",x"c0",x"98"),
  1603 => (x"48",x"66",x"c4",x"58"),
  1604 => (x"a6",x"cc",x"80",x"c4"),
  1605 => (x"bf",x"66",x"c8",x"58"),
  1606 => (x"66",x"e4",x"c0",x"4c"),
  1607 => (x"a8",x"66",x"cc",x"48"),
  1608 => (x"87",x"c5",x"c0",x"02"),
  1609 => (x"c2",x"c0",x"7e",x"c0"),
  1610 => (x"6e",x"7e",x"c1",x"87"),
  1611 => (x"1e",x"e0",x"c0",x"1e"),
  1612 => (x"d5",x"ff",x"49",x"74"),
  1613 => (x"86",x"c8",x"87",x"f6"),
  1614 => (x"b7",x"c0",x"4d",x"70"),
  1615 => (x"d4",x"c1",x"06",x"ad"),
  1616 => (x"c8",x"84",x"75",x"87"),
  1617 => (x"c0",x"49",x"bf",x"66"),
  1618 => (x"89",x"74",x"81",x"e0"),
  1619 => (x"fc",x"c9",x"c1",x"4b"),
  1620 => (x"de",x"fe",x"71",x"4a"),
  1621 => (x"84",x"c2",x"87",x"ea"),
  1622 => (x"e8",x"c0",x"7e",x"74"),
  1623 => (x"80",x"c1",x"48",x"66"),
  1624 => (x"58",x"a6",x"ec",x"c0"),
  1625 => (x"49",x"66",x"f0",x"c0"),
  1626 => (x"a9",x"70",x"81",x"c1"),
  1627 => (x"87",x"c5",x"c0",x"02"),
  1628 => (x"c2",x"c0",x"4c",x"c0"),
  1629 => (x"74",x"4c",x"c1",x"87"),
  1630 => (x"bf",x"66",x"cc",x"1e"),
  1631 => (x"81",x"e0",x"c0",x"49"),
  1632 => (x"71",x"89",x"66",x"c4"),
  1633 => (x"49",x"66",x"c8",x"1e"),
  1634 => (x"87",x"e0",x"d4",x"ff"),
  1635 => (x"b7",x"c0",x"86",x"c8"),
  1636 => (x"c5",x"ff",x"01",x"a8"),
  1637 => (x"66",x"e8",x"c0",x"87"),
  1638 => (x"87",x"d3",x"c0",x"02"),
  1639 => (x"c9",x"49",x"66",x"c4"),
  1640 => (x"66",x"e8",x"c0",x"81"),
  1641 => (x"48",x"66",x"c4",x"51"),
  1642 => (x"78",x"fe",x"d5",x"c1"),
  1643 => (x"c4",x"87",x"ce",x"c0"),
  1644 => (x"81",x"c9",x"49",x"66"),
  1645 => (x"66",x"c4",x"51",x"c2"),
  1646 => (x"fc",x"d7",x"c1",x"48"),
  1647 => (x"48",x"66",x"d4",x"78"),
  1648 => (x"04",x"a8",x"66",x"d8"),
  1649 => (x"d4",x"87",x"cb",x"c0"),
  1650 => (x"80",x"c1",x"48",x"66"),
  1651 => (x"c0",x"58",x"a6",x"d8"),
  1652 => (x"66",x"d8",x"87",x"d1"),
  1653 => (x"dc",x"88",x"c1",x"48"),
  1654 => (x"c6",x"c0",x"58",x"a6"),
  1655 => (x"f7",x"d2",x"ff",x"87"),
  1656 => (x"cc",x"4d",x"70",x"87"),
  1657 => (x"78",x"c0",x"48",x"a6"),
  1658 => (x"ff",x"87",x"c6",x"c0"),
  1659 => (x"70",x"87",x"e9",x"d2"),
  1660 => (x"66",x"e0",x"c0",x"4d"),
  1661 => (x"c0",x"80",x"c1",x"48"),
  1662 => (x"75",x"58",x"a6",x"e4"),
  1663 => (x"cb",x"c0",x"02",x"9d"),
  1664 => (x"48",x"66",x"d4",x"87"),
  1665 => (x"a8",x"66",x"cc",x"c1"),
  1666 => (x"87",x"da",x"f4",x"04"),
  1667 => (x"c7",x"48",x"66",x"d4"),
  1668 => (x"e1",x"c0",x"03",x"a8"),
  1669 => (x"4c",x"66",x"d4",x"87"),
  1670 => (x"48",x"c4",x"f3",x"c2"),
  1671 => (x"49",x"74",x"78",x"c0"),
  1672 => (x"c4",x"c1",x"91",x"cc"),
  1673 => (x"a1",x"c4",x"81",x"66"),
  1674 => (x"c0",x"4a",x"6a",x"4a"),
  1675 => (x"84",x"c1",x"79",x"52"),
  1676 => (x"ff",x"04",x"ac",x"c7"),
  1677 => (x"e4",x"c0",x"87",x"e2"),
  1678 => (x"e2",x"c0",x"02",x"66"),
  1679 => (x"66",x"c4",x"c1",x"87"),
  1680 => (x"81",x"d4",x"c1",x"49"),
  1681 => (x"4a",x"66",x"c4",x"c1"),
  1682 => (x"c0",x"82",x"dc",x"c1"),
  1683 => (x"f0",x"d4",x"c1",x"52"),
  1684 => (x"66",x"c4",x"c1",x"79"),
  1685 => (x"81",x"d8",x"c1",x"49"),
  1686 => (x"79",x"c0",x"ca",x"c1"),
  1687 => (x"c1",x"87",x"d6",x"c0"),
  1688 => (x"c1",x"49",x"66",x"c4"),
  1689 => (x"c4",x"c1",x"81",x"d4"),
  1690 => (x"d8",x"c1",x"4a",x"66"),
  1691 => (x"c8",x"ca",x"c1",x"82"),
  1692 => (x"e7",x"d4",x"c1",x"7a"),
  1693 => (x"66",x"c4",x"c1",x"79"),
  1694 => (x"81",x"e0",x"c1",x"49"),
  1695 => (x"79",x"ce",x"d8",x"c1"),
  1696 => (x"87",x"cb",x"d0",x"ff"),
  1697 => (x"ff",x"48",x"66",x"d0"),
  1698 => (x"4d",x"26",x"8e",x"cc"),
  1699 => (x"4b",x"26",x"4c",x"26"),
  1700 => (x"c7",x"1e",x"4f",x"26"),
  1701 => (x"c0",x"f3",x"c2",x"1e"),
  1702 => (x"ed",x"c1",x"1e",x"bf"),
  1703 => (x"f1",x"c2",x"1e",x"cc"),
  1704 => (x"49",x"bf",x"97",x"f0"),
  1705 => (x"c1",x"87",x"f9",x"ee"),
  1706 => (x"c0",x"49",x"cc",x"ed"),
  1707 => (x"f4",x"87",x"ff",x"e1"),
  1708 => (x"1e",x"4f",x"26",x"8e"),
  1709 => (x"48",x"c0",x"ed",x"c1"),
  1710 => (x"e3",x"c2",x"50",x"c0"),
  1711 => (x"ff",x"49",x"bf",x"e0"),
  1712 => (x"c0",x"87",x"c3",x"d5"),
  1713 => (x"1e",x"4f",x"26",x"48"),
  1714 => (x"cd",x"c7",x"1e",x"73"),
  1715 => (x"cc",x"f3",x"c2",x"87"),
  1716 => (x"ff",x"50",x"c0",x"48"),
  1717 => (x"ff",x"c3",x"48",x"d4"),
  1718 => (x"d0",x"ca",x"c1",x"78"),
  1719 => (x"c6",x"d7",x"fe",x"49"),
  1720 => (x"db",x"e2",x"fe",x"87"),
  1721 => (x"02",x"98",x"70",x"87"),
  1722 => (x"eb",x"fe",x"87",x"cd"),
  1723 => (x"98",x"70",x"87",x"f9"),
  1724 => (x"c1",x"87",x"c4",x"02"),
  1725 => (x"c0",x"87",x"c2",x"4a"),
  1726 => (x"02",x"9a",x"72",x"4a"),
  1727 => (x"ca",x"c1",x"87",x"c8"),
  1728 => (x"d6",x"fe",x"49",x"dc"),
  1729 => (x"f3",x"c2",x"87",x"e1"),
  1730 => (x"78",x"c0",x"48",x"c0"),
  1731 => (x"48",x"f0",x"f1",x"c2"),
  1732 => (x"fd",x"49",x"50",x"c0"),
  1733 => (x"da",x"fe",x"87",x"fc"),
  1734 => (x"9b",x"4b",x"70",x"87"),
  1735 => (x"c1",x"87",x"cf",x"02"),
  1736 => (x"c7",x"5b",x"e8",x"ee"),
  1737 => (x"87",x"f8",x"de",x"49"),
  1738 => (x"e0",x"c0",x"49",x"c1"),
  1739 => (x"f2",x"c2",x"87",x"d3"),
  1740 => (x"d9",x"e1",x"c0",x"87"),
  1741 => (x"f8",x"ef",x"c0",x"87"),
  1742 => (x"87",x"f5",x"ff",x"87"),
  1743 => (x"4f",x"26",x"4b",x"26"),
  1744 => (x"00",x"00",x"00",x"00"),
  1745 => (x"00",x"00",x"00",x"00"),
  1746 => (x"00",x"00",x"00",x"01"),
  1747 => (x"00",x"00",x"11",x"da"),
  1748 => (x"00",x"00",x"2c",x"d8"),
  1749 => (x"b4",x"00",x"00",x"00"),
  1750 => (x"00",x"00",x"11",x"da"),
  1751 => (x"00",x"00",x"2c",x"f6"),
  1752 => (x"b4",x"00",x"00",x"00"),
  1753 => (x"00",x"00",x"11",x"da"),
  1754 => (x"00",x"00",x"2d",x"14"),
  1755 => (x"b4",x"00",x"00",x"00"),
  1756 => (x"00",x"00",x"11",x"da"),
  1757 => (x"00",x"00",x"2d",x"32"),
  1758 => (x"b4",x"00",x"00",x"00"),
  1759 => (x"00",x"00",x"11",x"da"),
  1760 => (x"00",x"00",x"2d",x"50"),
  1761 => (x"b4",x"00",x"00",x"00"),
  1762 => (x"00",x"00",x"11",x"da"),
  1763 => (x"00",x"00",x"2d",x"6e"),
  1764 => (x"b4",x"00",x"00",x"00"),
  1765 => (x"00",x"00",x"11",x"da"),
  1766 => (x"00",x"00",x"2d",x"8c"),
  1767 => (x"b4",x"00",x"00",x"00"),
  1768 => (x"00",x"00",x"15",x"30"),
  1769 => (x"00",x"00",x"00",x"00"),
  1770 => (x"b4",x"00",x"00",x"00"),
  1771 => (x"00",x"00",x"12",x"d4"),
  1772 => (x"00",x"00",x"00",x"00"),
  1773 => (x"b4",x"00",x"00",x"00"),
  1774 => (x"00",x"00",x"12",x"a0"),
  1775 => (x"db",x"86",x"fc",x"1e"),
  1776 => (x"fc",x"7e",x"70",x"87"),
  1777 => (x"1e",x"4f",x"26",x"8e"),
  1778 => (x"c0",x"48",x"f0",x"fe"),
  1779 => (x"79",x"09",x"cd",x"78"),
  1780 => (x"1e",x"4f",x"26",x"09"),
  1781 => (x"49",x"fc",x"ee",x"c1"),
  1782 => (x"4f",x"26",x"87",x"ed"),
  1783 => (x"bf",x"f0",x"fe",x"1e"),
  1784 => (x"1e",x"4f",x"26",x"48"),
  1785 => (x"c1",x"48",x"f0",x"fe"),
  1786 => (x"1e",x"4f",x"26",x"78"),
  1787 => (x"c0",x"48",x"f0",x"fe"),
  1788 => (x"1e",x"4f",x"26",x"78"),
  1789 => (x"52",x"c0",x"4a",x"71"),
  1790 => (x"0e",x"4f",x"26",x"51"),
  1791 => (x"5d",x"5c",x"5b",x"5e"),
  1792 => (x"71",x"86",x"f4",x"0e"),
  1793 => (x"7e",x"6d",x"97",x"4d"),
  1794 => (x"97",x"4c",x"a5",x"c1"),
  1795 => (x"a6",x"c8",x"48",x"6c"),
  1796 => (x"c4",x"48",x"6e",x"58"),
  1797 => (x"c5",x"05",x"a8",x"66"),
  1798 => (x"c0",x"48",x"ff",x"87"),
  1799 => (x"ca",x"ff",x"87",x"e6"),
  1800 => (x"49",x"a5",x"c2",x"87"),
  1801 => (x"71",x"4b",x"6c",x"97"),
  1802 => (x"6b",x"97",x"4b",x"a3"),
  1803 => (x"7e",x"6c",x"97",x"4b"),
  1804 => (x"80",x"c1",x"48",x"6e"),
  1805 => (x"c7",x"58",x"a6",x"c8"),
  1806 => (x"58",x"a6",x"cc",x"98"),
  1807 => (x"fe",x"7c",x"97",x"70"),
  1808 => (x"48",x"73",x"87",x"e1"),
  1809 => (x"4d",x"26",x"8e",x"f4"),
  1810 => (x"4b",x"26",x"4c",x"26"),
  1811 => (x"73",x"1e",x"4f",x"26"),
  1812 => (x"fe",x"86",x"f4",x"1e"),
  1813 => (x"bf",x"e0",x"87",x"d5"),
  1814 => (x"e0",x"c0",x"49",x"4b"),
  1815 => (x"c0",x"02",x"99",x"c0"),
  1816 => (x"4a",x"73",x"87",x"ea"),
  1817 => (x"c2",x"9a",x"ff",x"c3"),
  1818 => (x"bf",x"97",x"c0",x"f7"),
  1819 => (x"c2",x"f7",x"c2",x"49"),
  1820 => (x"c2",x"51",x"72",x"81"),
  1821 => (x"bf",x"97",x"c0",x"f7"),
  1822 => (x"c1",x"48",x"6e",x"7e"),
  1823 => (x"58",x"a6",x"c8",x"80"),
  1824 => (x"a6",x"cc",x"98",x"c7"),
  1825 => (x"c0",x"f7",x"c2",x"58"),
  1826 => (x"50",x"66",x"c8",x"48"),
  1827 => (x"70",x"87",x"cd",x"fd"),
  1828 => (x"87",x"cf",x"fd",x"7e"),
  1829 => (x"4b",x"26",x"8e",x"f4"),
  1830 => (x"c2",x"1e",x"4f",x"26"),
  1831 => (x"fd",x"49",x"c0",x"f7"),
  1832 => (x"f1",x"c1",x"87",x"d1"),
  1833 => (x"de",x"fc",x"49",x"ce"),
  1834 => (x"87",x"e8",x"c4",x"87"),
  1835 => (x"5e",x"0e",x"4f",x"26"),
  1836 => (x"0e",x"5d",x"5c",x"5b"),
  1837 => (x"7e",x"71",x"86",x"fc"),
  1838 => (x"c2",x"4d",x"d4",x"ff"),
  1839 => (x"fc",x"49",x"c0",x"f7"),
  1840 => (x"4b",x"70",x"87",x"f9"),
  1841 => (x"04",x"ab",x"b7",x"c0"),
  1842 => (x"c3",x"87",x"f5",x"c2"),
  1843 => (x"c9",x"05",x"ab",x"f0"),
  1844 => (x"cc",x"f6",x"c1",x"87"),
  1845 => (x"c2",x"78",x"c1",x"48"),
  1846 => (x"e0",x"c3",x"87",x"d6"),
  1847 => (x"87",x"c9",x"05",x"ab"),
  1848 => (x"48",x"d0",x"f6",x"c1"),
  1849 => (x"c7",x"c2",x"78",x"c1"),
  1850 => (x"d0",x"f6",x"c1",x"87"),
  1851 => (x"87",x"c6",x"02",x"bf"),
  1852 => (x"4c",x"a3",x"c0",x"c2"),
  1853 => (x"4c",x"73",x"87",x"c2"),
  1854 => (x"bf",x"cc",x"f6",x"c1"),
  1855 => (x"87",x"e0",x"c0",x"02"),
  1856 => (x"b7",x"c4",x"49",x"74"),
  1857 => (x"f6",x"c1",x"91",x"29"),
  1858 => (x"4a",x"74",x"81",x"d4"),
  1859 => (x"92",x"c2",x"9a",x"cf"),
  1860 => (x"30",x"72",x"48",x"c1"),
  1861 => (x"ba",x"ff",x"4a",x"70"),
  1862 => (x"98",x"69",x"48",x"72"),
  1863 => (x"87",x"db",x"79",x"70"),
  1864 => (x"b7",x"c4",x"49",x"74"),
  1865 => (x"f6",x"c1",x"91",x"29"),
  1866 => (x"4a",x"74",x"81",x"d4"),
  1867 => (x"92",x"c2",x"9a",x"cf"),
  1868 => (x"30",x"72",x"48",x"c3"),
  1869 => (x"69",x"48",x"4a",x"70"),
  1870 => (x"6e",x"79",x"70",x"b0"),
  1871 => (x"87",x"e4",x"c0",x"05"),
  1872 => (x"c8",x"48",x"d0",x"ff"),
  1873 => (x"7d",x"c5",x"78",x"e1"),
  1874 => (x"bf",x"d0",x"f6",x"c1"),
  1875 => (x"c3",x"87",x"c3",x"02"),
  1876 => (x"f6",x"c1",x"7d",x"e0"),
  1877 => (x"c3",x"02",x"bf",x"cc"),
  1878 => (x"7d",x"f0",x"c3",x"87"),
  1879 => (x"d0",x"ff",x"7d",x"73"),
  1880 => (x"78",x"e0",x"c0",x"48"),
  1881 => (x"48",x"d0",x"f6",x"c1"),
  1882 => (x"f6",x"c1",x"78",x"c0"),
  1883 => (x"78",x"c0",x"48",x"cc"),
  1884 => (x"49",x"c0",x"f7",x"c2"),
  1885 => (x"70",x"87",x"c4",x"fa"),
  1886 => (x"ab",x"b7",x"c0",x"4b"),
  1887 => (x"87",x"cb",x"fd",x"03"),
  1888 => (x"8e",x"fc",x"48",x"c0"),
  1889 => (x"4c",x"26",x"4d",x"26"),
  1890 => (x"4f",x"26",x"4b",x"26"),
  1891 => (x"00",x"00",x"00",x"00"),
  1892 => (x"00",x"00",x"00",x"00"),
  1893 => (x"00",x"00",x"00",x"00"),
  1894 => (x"34",x"34",x"34",x"34"),
  1895 => (x"34",x"34",x"34",x"34"),
  1896 => (x"34",x"34",x"34",x"34"),
  1897 => (x"34",x"34",x"34",x"34"),
  1898 => (x"34",x"34",x"34",x"34"),
  1899 => (x"34",x"34",x"34",x"34"),
  1900 => (x"34",x"34",x"34",x"34"),
  1901 => (x"34",x"34",x"34",x"34"),
  1902 => (x"34",x"34",x"34",x"34"),
  1903 => (x"34",x"34",x"34",x"34"),
  1904 => (x"34",x"34",x"34",x"34"),
  1905 => (x"34",x"34",x"34",x"34"),
  1906 => (x"34",x"34",x"34",x"34"),
  1907 => (x"34",x"34",x"34",x"34"),
  1908 => (x"34",x"34",x"34",x"34"),
  1909 => (x"72",x"4a",x"c0",x"1e"),
  1910 => (x"c1",x"91",x"c4",x"49"),
  1911 => (x"c0",x"81",x"d4",x"f6"),
  1912 => (x"d0",x"82",x"c1",x"79"),
  1913 => (x"ee",x"04",x"aa",x"b7"),
  1914 => (x"0e",x"4f",x"26",x"87"),
  1915 => (x"5d",x"5c",x"5b",x"5e"),
  1916 => (x"f7",x"4d",x"71",x"0e"),
  1917 => (x"4a",x"75",x"87",x"f5"),
  1918 => (x"92",x"2a",x"b7",x"c4"),
  1919 => (x"82",x"d4",x"f6",x"c1"),
  1920 => (x"9c",x"cf",x"4c",x"75"),
  1921 => (x"49",x"6a",x"94",x"c2"),
  1922 => (x"c3",x"2b",x"74",x"4b"),
  1923 => (x"74",x"48",x"c2",x"9b"),
  1924 => (x"ff",x"4c",x"70",x"30"),
  1925 => (x"71",x"48",x"74",x"bc"),
  1926 => (x"f7",x"7a",x"70",x"98"),
  1927 => (x"48",x"73",x"87",x"c5"),
  1928 => (x"4c",x"26",x"4d",x"26"),
  1929 => (x"4f",x"26",x"4b",x"26"),
  1930 => (x"48",x"d0",x"ff",x"1e"),
  1931 => (x"71",x"78",x"e1",x"c8"),
  1932 => (x"08",x"d4",x"ff",x"48"),
  1933 => (x"1e",x"4f",x"26",x"78"),
  1934 => (x"c8",x"48",x"d0",x"ff"),
  1935 => (x"48",x"71",x"78",x"e1"),
  1936 => (x"78",x"08",x"d4",x"ff"),
  1937 => (x"ff",x"48",x"66",x"c4"),
  1938 => (x"26",x"78",x"08",x"d4"),
  1939 => (x"4a",x"71",x"1e",x"4f"),
  1940 => (x"1e",x"49",x"66",x"c4"),
  1941 => (x"de",x"ff",x"49",x"72"),
  1942 => (x"48",x"d0",x"ff",x"87"),
  1943 => (x"fc",x"78",x"e0",x"c0"),
  1944 => (x"1e",x"4f",x"26",x"8e"),
  1945 => (x"4a",x"71",x"1e",x"73"),
  1946 => (x"ab",x"b7",x"c2",x"4b"),
  1947 => (x"a3",x"87",x"c8",x"03"),
  1948 => (x"ff",x"c3",x"4a",x"49"),
  1949 => (x"ce",x"87",x"c7",x"9a"),
  1950 => (x"c3",x"4a",x"49",x"a3"),
  1951 => (x"66",x"c8",x"9a",x"ff"),
  1952 => (x"49",x"72",x"1e",x"49"),
  1953 => (x"fc",x"87",x"c6",x"ff"),
  1954 => (x"26",x"4b",x"26",x"8e"),
  1955 => (x"d0",x"ff",x"1e",x"4f"),
  1956 => (x"78",x"c9",x"c8",x"48"),
  1957 => (x"d4",x"ff",x"48",x"71"),
  1958 => (x"4f",x"26",x"78",x"08"),
  1959 => (x"49",x"4a",x"71",x"1e"),
  1960 => (x"d0",x"ff",x"87",x"eb"),
  1961 => (x"26",x"78",x"c8",x"48"),
  1962 => (x"1e",x"73",x"1e",x"4f"),
  1963 => (x"f7",x"c2",x"4b",x"71"),
  1964 => (x"c3",x"02",x"bf",x"d8"),
  1965 => (x"87",x"eb",x"c2",x"87"),
  1966 => (x"c8",x"48",x"d0",x"ff"),
  1967 => (x"48",x"73",x"78",x"c9"),
  1968 => (x"ff",x"b0",x"e0",x"c0"),
  1969 => (x"c2",x"78",x"08",x"d4"),
  1970 => (x"c0",x"48",x"cc",x"f7"),
  1971 => (x"02",x"66",x"c8",x"78"),
  1972 => (x"ff",x"c3",x"87",x"c5"),
  1973 => (x"c0",x"87",x"c2",x"49"),
  1974 => (x"d4",x"f7",x"c2",x"49"),
  1975 => (x"02",x"66",x"cc",x"59"),
  1976 => (x"d5",x"c5",x"87",x"c6"),
  1977 => (x"87",x"c4",x"4a",x"d5"),
  1978 => (x"4a",x"ff",x"ff",x"cf"),
  1979 => (x"5a",x"d8",x"f7",x"c2"),
  1980 => (x"48",x"d8",x"f7",x"c2"),
  1981 => (x"4b",x"26",x"78",x"c1"),
  1982 => (x"5e",x"0e",x"4f",x"26"),
  1983 => (x"0e",x"5d",x"5c",x"5b"),
  1984 => (x"f7",x"c2",x"4d",x"71"),
  1985 => (x"75",x"4b",x"bf",x"d4"),
  1986 => (x"87",x"cb",x"02",x"9d"),
  1987 => (x"c1",x"91",x"c8",x"49"),
  1988 => (x"71",x"4a",x"e0",x"fa"),
  1989 => (x"c1",x"87",x"c4",x"82"),
  1990 => (x"c0",x"4a",x"e0",x"fe"),
  1991 => (x"73",x"49",x"12",x"4c"),
  1992 => (x"d0",x"f7",x"c2",x"99"),
  1993 => (x"b8",x"71",x"48",x"bf"),
  1994 => (x"78",x"08",x"d4",x"ff"),
  1995 => (x"84",x"2b",x"b7",x"c1"),
  1996 => (x"04",x"ac",x"b7",x"c8"),
  1997 => (x"f7",x"c2",x"87",x"e7"),
  1998 => (x"c8",x"48",x"bf",x"cc"),
  1999 => (x"d0",x"f7",x"c2",x"80"),
  2000 => (x"26",x"4d",x"26",x"58"),
  2001 => (x"26",x"4b",x"26",x"4c"),
  2002 => (x"1e",x"73",x"1e",x"4f"),
  2003 => (x"4a",x"13",x"4b",x"71"),
  2004 => (x"87",x"cb",x"02",x"9a"),
  2005 => (x"e1",x"fe",x"49",x"72"),
  2006 => (x"9a",x"4a",x"13",x"87"),
  2007 => (x"26",x"87",x"f5",x"05"),
  2008 => (x"1e",x"4f",x"26",x"4b"),
  2009 => (x"bf",x"cc",x"f7",x"c2"),
  2010 => (x"cc",x"f7",x"c2",x"49"),
  2011 => (x"78",x"a1",x"c1",x"48"),
  2012 => (x"a9",x"b7",x"c0",x"c4"),
  2013 => (x"ff",x"87",x"db",x"03"),
  2014 => (x"f7",x"c2",x"48",x"d4"),
  2015 => (x"c2",x"78",x"bf",x"d0"),
  2016 => (x"49",x"bf",x"cc",x"f7"),
  2017 => (x"48",x"cc",x"f7",x"c2"),
  2018 => (x"c4",x"78",x"a1",x"c1"),
  2019 => (x"04",x"a9",x"b7",x"c0"),
  2020 => (x"d0",x"ff",x"87",x"e5"),
  2021 => (x"c2",x"78",x"c8",x"48"),
  2022 => (x"c0",x"48",x"d8",x"f7"),
  2023 => (x"00",x"4f",x"26",x"78"),
  2024 => (x"00",x"00",x"00",x"00"),
  2025 => (x"00",x"00",x"00",x"00"),
  2026 => (x"5f",x"00",x"00",x"00"),
  2027 => (x"00",x"00",x"00",x"5f"),
  2028 => (x"00",x"03",x"03",x"00"),
  2029 => (x"00",x"00",x"03",x"03"),
  2030 => (x"14",x"7f",x"7f",x"14"),
  2031 => (x"00",x"14",x"7f",x"7f"),
  2032 => (x"6b",x"2e",x"24",x"00"),
  2033 => (x"00",x"12",x"3a",x"6b"),
  2034 => (x"18",x"36",x"6a",x"4c"),
  2035 => (x"00",x"32",x"56",x"6c"),
  2036 => (x"59",x"4f",x"7e",x"30"),
  2037 => (x"40",x"68",x"3a",x"77"),
  2038 => (x"07",x"04",x"00",x"00"),
  2039 => (x"00",x"00",x"00",x"03"),
  2040 => (x"3e",x"1c",x"00",x"00"),
  2041 => (x"00",x"00",x"41",x"63"),
  2042 => (x"63",x"41",x"00",x"00"),
  2043 => (x"00",x"00",x"1c",x"3e"),
  2044 => (x"1c",x"3e",x"2a",x"08"),
  2045 => (x"08",x"2a",x"3e",x"1c"),
  2046 => (x"3e",x"08",x"08",x"00"),
  2047 => (x"00",x"08",x"08",x"3e"),
  2048 => (x"e0",x"80",x"00",x"00"),
  2049 => (x"00",x"00",x"00",x"60"),
  2050 => (x"08",x"08",x"08",x"00"),
  2051 => (x"00",x"08",x"08",x"08"),
  2052 => (x"60",x"00",x"00",x"00"),
  2053 => (x"00",x"00",x"00",x"60"),
  2054 => (x"18",x"30",x"60",x"40"),
  2055 => (x"01",x"03",x"06",x"0c"),
  2056 => (x"59",x"7f",x"3e",x"00"),
  2057 => (x"00",x"3e",x"7f",x"4d"),
  2058 => (x"7f",x"06",x"04",x"00"),
  2059 => (x"00",x"00",x"00",x"7f"),
  2060 => (x"71",x"63",x"42",x"00"),
  2061 => (x"00",x"46",x"4f",x"59"),
  2062 => (x"49",x"63",x"22",x"00"),
  2063 => (x"00",x"36",x"7f",x"49"),
  2064 => (x"13",x"16",x"1c",x"18"),
  2065 => (x"00",x"10",x"7f",x"7f"),
  2066 => (x"45",x"67",x"27",x"00"),
  2067 => (x"00",x"39",x"7d",x"45"),
  2068 => (x"4b",x"7e",x"3c",x"00"),
  2069 => (x"00",x"30",x"79",x"49"),
  2070 => (x"71",x"01",x"01",x"00"),
  2071 => (x"00",x"07",x"0f",x"79"),
  2072 => (x"49",x"7f",x"36",x"00"),
  2073 => (x"00",x"36",x"7f",x"49"),
  2074 => (x"49",x"4f",x"06",x"00"),
  2075 => (x"00",x"1e",x"3f",x"69"),
  2076 => (x"66",x"00",x"00",x"00"),
  2077 => (x"00",x"00",x"00",x"66"),
  2078 => (x"e6",x"80",x"00",x"00"),
  2079 => (x"00",x"00",x"00",x"66"),
  2080 => (x"14",x"08",x"08",x"00"),
  2081 => (x"00",x"22",x"22",x"14"),
  2082 => (x"14",x"14",x"14",x"00"),
  2083 => (x"00",x"14",x"14",x"14"),
  2084 => (x"14",x"22",x"22",x"00"),
  2085 => (x"00",x"08",x"08",x"14"),
  2086 => (x"51",x"03",x"02",x"00"),
  2087 => (x"00",x"06",x"0f",x"59"),
  2088 => (x"5d",x"41",x"7f",x"3e"),
  2089 => (x"00",x"1e",x"1f",x"55"),
  2090 => (x"09",x"7f",x"7e",x"00"),
  2091 => (x"00",x"7e",x"7f",x"09"),
  2092 => (x"49",x"7f",x"7f",x"00"),
  2093 => (x"00",x"36",x"7f",x"49"),
  2094 => (x"63",x"3e",x"1c",x"00"),
  2095 => (x"00",x"41",x"41",x"41"),
  2096 => (x"41",x"7f",x"7f",x"00"),
  2097 => (x"00",x"1c",x"3e",x"63"),
  2098 => (x"49",x"7f",x"7f",x"00"),
  2099 => (x"00",x"41",x"41",x"49"),
  2100 => (x"09",x"7f",x"7f",x"00"),
  2101 => (x"00",x"01",x"01",x"09"),
  2102 => (x"41",x"7f",x"3e",x"00"),
  2103 => (x"00",x"7a",x"7b",x"49"),
  2104 => (x"08",x"7f",x"7f",x"00"),
  2105 => (x"00",x"7f",x"7f",x"08"),
  2106 => (x"7f",x"41",x"00",x"00"),
  2107 => (x"00",x"00",x"41",x"7f"),
  2108 => (x"40",x"60",x"20",x"00"),
  2109 => (x"00",x"3f",x"7f",x"40"),
  2110 => (x"1c",x"08",x"7f",x"7f"),
  2111 => (x"00",x"41",x"63",x"36"),
  2112 => (x"40",x"7f",x"7f",x"00"),
  2113 => (x"00",x"40",x"40",x"40"),
  2114 => (x"0c",x"06",x"7f",x"7f"),
  2115 => (x"00",x"7f",x"7f",x"06"),
  2116 => (x"0c",x"06",x"7f",x"7f"),
  2117 => (x"00",x"7f",x"7f",x"18"),
  2118 => (x"41",x"7f",x"3e",x"00"),
  2119 => (x"00",x"3e",x"7f",x"41"),
  2120 => (x"09",x"7f",x"7f",x"00"),
  2121 => (x"00",x"06",x"0f",x"09"),
  2122 => (x"61",x"41",x"7f",x"3e"),
  2123 => (x"00",x"40",x"7e",x"7f"),
  2124 => (x"09",x"7f",x"7f",x"00"),
  2125 => (x"00",x"66",x"7f",x"19"),
  2126 => (x"4d",x"6f",x"26",x"00"),
  2127 => (x"00",x"32",x"7b",x"59"),
  2128 => (x"7f",x"01",x"01",x"00"),
  2129 => (x"00",x"01",x"01",x"7f"),
  2130 => (x"40",x"7f",x"3f",x"00"),
  2131 => (x"00",x"3f",x"7f",x"40"),
  2132 => (x"70",x"3f",x"0f",x"00"),
  2133 => (x"00",x"0f",x"3f",x"70"),
  2134 => (x"18",x"30",x"7f",x"7f"),
  2135 => (x"00",x"7f",x"7f",x"30"),
  2136 => (x"1c",x"36",x"63",x"41"),
  2137 => (x"41",x"63",x"36",x"1c"),
  2138 => (x"7c",x"06",x"03",x"01"),
  2139 => (x"01",x"03",x"06",x"7c"),
  2140 => (x"4d",x"59",x"71",x"61"),
  2141 => (x"00",x"41",x"43",x"47"),
  2142 => (x"7f",x"7f",x"00",x"00"),
  2143 => (x"00",x"00",x"41",x"41"),
  2144 => (x"0c",x"06",x"03",x"01"),
  2145 => (x"40",x"60",x"30",x"18"),
  2146 => (x"41",x"41",x"00",x"00"),
  2147 => (x"00",x"00",x"7f",x"7f"),
  2148 => (x"03",x"06",x"0c",x"08"),
  2149 => (x"00",x"08",x"0c",x"06"),
  2150 => (x"80",x"80",x"80",x"80"),
  2151 => (x"00",x"80",x"80",x"80"),
  2152 => (x"03",x"00",x"00",x"00"),
  2153 => (x"00",x"00",x"04",x"07"),
  2154 => (x"54",x"74",x"20",x"00"),
  2155 => (x"00",x"78",x"7c",x"54"),
  2156 => (x"44",x"7f",x"7f",x"00"),
  2157 => (x"00",x"38",x"7c",x"44"),
  2158 => (x"44",x"7c",x"38",x"00"),
  2159 => (x"00",x"00",x"44",x"44"),
  2160 => (x"44",x"7c",x"38",x"00"),
  2161 => (x"00",x"7f",x"7f",x"44"),
  2162 => (x"54",x"7c",x"38",x"00"),
  2163 => (x"00",x"18",x"5c",x"54"),
  2164 => (x"7f",x"7e",x"04",x"00"),
  2165 => (x"00",x"00",x"05",x"05"),
  2166 => (x"a4",x"bc",x"18",x"00"),
  2167 => (x"00",x"7c",x"fc",x"a4"),
  2168 => (x"04",x"7f",x"7f",x"00"),
  2169 => (x"00",x"78",x"7c",x"04"),
  2170 => (x"3d",x"00",x"00",x"00"),
  2171 => (x"00",x"00",x"40",x"7d"),
  2172 => (x"80",x"80",x"80",x"00"),
  2173 => (x"00",x"00",x"7d",x"fd"),
  2174 => (x"10",x"7f",x"7f",x"00"),
  2175 => (x"00",x"44",x"6c",x"38"),
  2176 => (x"3f",x"00",x"00",x"00"),
  2177 => (x"00",x"00",x"40",x"7f"),
  2178 => (x"18",x"0c",x"7c",x"7c"),
  2179 => (x"00",x"78",x"7c",x"0c"),
  2180 => (x"04",x"7c",x"7c",x"00"),
  2181 => (x"00",x"78",x"7c",x"04"),
  2182 => (x"44",x"7c",x"38",x"00"),
  2183 => (x"00",x"38",x"7c",x"44"),
  2184 => (x"24",x"fc",x"fc",x"00"),
  2185 => (x"00",x"18",x"3c",x"24"),
  2186 => (x"24",x"3c",x"18",x"00"),
  2187 => (x"00",x"fc",x"fc",x"24"),
  2188 => (x"04",x"7c",x"7c",x"00"),
  2189 => (x"00",x"08",x"0c",x"04"),
  2190 => (x"54",x"5c",x"48",x"00"),
  2191 => (x"00",x"20",x"74",x"54"),
  2192 => (x"7f",x"3f",x"04",x"00"),
  2193 => (x"00",x"00",x"44",x"44"),
  2194 => (x"40",x"7c",x"3c",x"00"),
  2195 => (x"00",x"7c",x"7c",x"40"),
  2196 => (x"60",x"3c",x"1c",x"00"),
  2197 => (x"00",x"1c",x"3c",x"60"),
  2198 => (x"30",x"60",x"7c",x"3c"),
  2199 => (x"00",x"3c",x"7c",x"60"),
  2200 => (x"10",x"38",x"6c",x"44"),
  2201 => (x"00",x"44",x"6c",x"38"),
  2202 => (x"e0",x"bc",x"1c",x"00"),
  2203 => (x"00",x"1c",x"3c",x"60"),
  2204 => (x"74",x"64",x"44",x"00"),
  2205 => (x"00",x"44",x"4c",x"5c"),
  2206 => (x"3e",x"08",x"08",x"00"),
  2207 => (x"00",x"41",x"41",x"77"),
  2208 => (x"7f",x"00",x"00",x"00"),
  2209 => (x"00",x"00",x"00",x"7f"),
  2210 => (x"77",x"41",x"41",x"00"),
  2211 => (x"00",x"08",x"08",x"3e"),
  2212 => (x"03",x"01",x"01",x"02"),
  2213 => (x"00",x"01",x"02",x"02"),
  2214 => (x"7f",x"7f",x"7f",x"7f"),
  2215 => (x"00",x"7f",x"7f",x"7f"),
  2216 => (x"1c",x"1c",x"08",x"08"),
  2217 => (x"7f",x"7f",x"3e",x"3e"),
  2218 => (x"3e",x"3e",x"7f",x"7f"),
  2219 => (x"08",x"08",x"1c",x"1c"),
  2220 => (x"7c",x"18",x"10",x"00"),
  2221 => (x"00",x"10",x"18",x"7c"),
  2222 => (x"7c",x"30",x"10",x"00"),
  2223 => (x"00",x"10",x"30",x"7c"),
  2224 => (x"60",x"60",x"30",x"10"),
  2225 => (x"00",x"06",x"1e",x"78"),
  2226 => (x"18",x"3c",x"66",x"42"),
  2227 => (x"00",x"42",x"66",x"3c"),
  2228 => (x"c2",x"6a",x"38",x"78"),
  2229 => (x"00",x"38",x"6c",x"c6"),
  2230 => (x"60",x"00",x"00",x"60"),
  2231 => (x"00",x"60",x"00",x"00"),
  2232 => (x"5c",x"5b",x"5e",x"0e"),
  2233 => (x"86",x"fc",x"0e",x"5d"),
  2234 => (x"f7",x"c2",x"7e",x"71"),
  2235 => (x"c0",x"4c",x"bf",x"e0"),
  2236 => (x"c4",x"1e",x"c0",x"4b"),
  2237 => (x"c4",x"02",x"ab",x"66"),
  2238 => (x"c2",x"4d",x"c0",x"87"),
  2239 => (x"75",x"4d",x"c1",x"87"),
  2240 => (x"ee",x"49",x"73",x"1e"),
  2241 => (x"86",x"c8",x"87",x"e3"),
  2242 => (x"ef",x"49",x"e0",x"c0"),
  2243 => (x"a4",x"c4",x"87",x"ec"),
  2244 => (x"f0",x"49",x"6a",x"4a"),
  2245 => (x"ca",x"f1",x"87",x"f3"),
  2246 => (x"c1",x"84",x"cc",x"87"),
  2247 => (x"ab",x"b7",x"c8",x"83"),
  2248 => (x"87",x"cd",x"ff",x"04"),
  2249 => (x"4d",x"26",x"8e",x"fc"),
  2250 => (x"4b",x"26",x"4c",x"26"),
  2251 => (x"71",x"1e",x"4f",x"26"),
  2252 => (x"e4",x"f7",x"c2",x"4a"),
  2253 => (x"e4",x"f7",x"c2",x"5a"),
  2254 => (x"49",x"78",x"c7",x"48"),
  2255 => (x"26",x"87",x"e1",x"fe"),
  2256 => (x"1e",x"73",x"1e",x"4f"),
  2257 => (x"0b",x"fc",x"4b",x"71"),
  2258 => (x"4a",x"73",x"0b",x"7b"),
  2259 => (x"c0",x"c1",x"9a",x"c1"),
  2260 => (x"c7",x"ed",x"49",x"a2"),
  2261 => (x"d8",x"da",x"c2",x"87"),
  2262 => (x"26",x"4b",x"26",x"5b"),
  2263 => (x"4a",x"71",x"1e",x"4f"),
  2264 => (x"72",x"1e",x"66",x"c4"),
  2265 => (x"87",x"fb",x"eb",x"49"),
  2266 => (x"4f",x"26",x"8e",x"fc"),
  2267 => (x"48",x"d4",x"ff",x"1e"),
  2268 => (x"ff",x"78",x"ff",x"c3"),
  2269 => (x"e1",x"c0",x"48",x"d0"),
  2270 => (x"48",x"d4",x"ff",x"78"),
  2271 => (x"48",x"71",x"78",x"c1"),
  2272 => (x"d4",x"ff",x"30",x"c4"),
  2273 => (x"d0",x"ff",x"78",x"08"),
  2274 => (x"78",x"e0",x"c0",x"48"),
  2275 => (x"5e",x"0e",x"4f",x"26"),
  2276 => (x"0e",x"5d",x"5c",x"5b"),
  2277 => (x"7e",x"c0",x"86",x"f4"),
  2278 => (x"ec",x"48",x"a6",x"c8"),
  2279 => (x"80",x"fc",x"78",x"bf"),
  2280 => (x"bf",x"e0",x"f7",x"c2"),
  2281 => (x"e8",x"f7",x"c2",x"78"),
  2282 => (x"bf",x"e8",x"4c",x"bf"),
  2283 => (x"d4",x"da",x"c2",x"4d"),
  2284 => (x"f9",x"e3",x"49",x"bf"),
  2285 => (x"e8",x"49",x"c7",x"87"),
  2286 => (x"49",x"70",x"87",x"f1"),
  2287 => (x"d0",x"05",x"99",x"c2"),
  2288 => (x"cc",x"da",x"c2",x"87"),
  2289 => (x"b9",x"ff",x"49",x"bf"),
  2290 => (x"c1",x"99",x"66",x"c8"),
  2291 => (x"f9",x"c1",x"02",x"99"),
  2292 => (x"49",x"e8",x"cf",x"87"),
  2293 => (x"70",x"87",x"c1",x"cb"),
  2294 => (x"e8",x"49",x"c7",x"4b"),
  2295 => (x"98",x"70",x"87",x"cd"),
  2296 => (x"c8",x"87",x"c9",x"05"),
  2297 => (x"99",x"c1",x"49",x"66"),
  2298 => (x"87",x"fe",x"c0",x"02"),
  2299 => (x"ec",x"48",x"a6",x"c8"),
  2300 => (x"f9",x"e2",x"78",x"bf"),
  2301 => (x"ca",x"49",x"73",x"87"),
  2302 => (x"98",x"70",x"87",x"ea"),
  2303 => (x"c2",x"87",x"d7",x"02"),
  2304 => (x"49",x"bf",x"c8",x"da"),
  2305 => (x"da",x"c2",x"b9",x"c1"),
  2306 => (x"fd",x"71",x"59",x"cc"),
  2307 => (x"e8",x"cf",x"87",x"de"),
  2308 => (x"87",x"c4",x"ca",x"49"),
  2309 => (x"49",x"c7",x"4b",x"70"),
  2310 => (x"70",x"87",x"d0",x"e7"),
  2311 => (x"cb",x"ff",x"05",x"98"),
  2312 => (x"49",x"66",x"c8",x"87"),
  2313 => (x"ff",x"05",x"99",x"c1"),
  2314 => (x"da",x"c2",x"87",x"c2"),
  2315 => (x"c1",x"4a",x"bf",x"d4"),
  2316 => (x"d8",x"da",x"c2",x"ba"),
  2317 => (x"7a",x"0a",x"fc",x"5a"),
  2318 => (x"c1",x"9a",x"c1",x"0a"),
  2319 => (x"e9",x"49",x"a2",x"c0"),
  2320 => (x"da",x"c1",x"87",x"da"),
  2321 => (x"87",x"e3",x"e6",x"49"),
  2322 => (x"da",x"c2",x"7e",x"c1"),
  2323 => (x"66",x"c8",x"48",x"cc"),
  2324 => (x"d4",x"da",x"c2",x"78"),
  2325 => (x"e9",x"c0",x"05",x"bf"),
  2326 => (x"c3",x"49",x"75",x"87"),
  2327 => (x"1e",x"71",x"99",x"ff"),
  2328 => (x"f8",x"fb",x"49",x"c0"),
  2329 => (x"c8",x"49",x"75",x"87"),
  2330 => (x"1e",x"71",x"29",x"b7"),
  2331 => (x"ec",x"fb",x"49",x"c1"),
  2332 => (x"c3",x"86",x"c8",x"87"),
  2333 => (x"f2",x"e5",x"49",x"fd"),
  2334 => (x"49",x"fa",x"c3",x"87"),
  2335 => (x"c7",x"87",x"ec",x"e5"),
  2336 => (x"49",x"75",x"87",x"f5"),
  2337 => (x"c8",x"99",x"ff",x"c3"),
  2338 => (x"b5",x"71",x"2d",x"b7"),
  2339 => (x"c0",x"02",x"9d",x"75"),
  2340 => (x"a6",x"c8",x"87",x"e4"),
  2341 => (x"bf",x"c8",x"ff",x"48"),
  2342 => (x"49",x"66",x"c8",x"78"),
  2343 => (x"bf",x"d0",x"da",x"c2"),
  2344 => (x"a9",x"e0",x"c2",x"89"),
  2345 => (x"87",x"c4",x"c0",x"03"),
  2346 => (x"87",x"d0",x"4d",x"c0"),
  2347 => (x"48",x"d0",x"da",x"c2"),
  2348 => (x"c0",x"78",x"66",x"c8"),
  2349 => (x"da",x"c2",x"87",x"c6"),
  2350 => (x"78",x"c0",x"48",x"d0"),
  2351 => (x"99",x"c8",x"49",x"75"),
  2352 => (x"87",x"ce",x"c0",x"05"),
  2353 => (x"e4",x"49",x"f5",x"c3"),
  2354 => (x"49",x"70",x"87",x"e1"),
  2355 => (x"c0",x"02",x"99",x"c2"),
  2356 => (x"f7",x"c2",x"87",x"e7"),
  2357 => (x"c0",x"02",x"bf",x"e4"),
  2358 => (x"c1",x"48",x"87",x"ca"),
  2359 => (x"e8",x"f7",x"c2",x"88"),
  2360 => (x"87",x"d3",x"c0",x"58"),
  2361 => (x"c1",x"48",x"66",x"c4"),
  2362 => (x"7e",x"70",x"80",x"e0"),
  2363 => (x"c0",x"02",x"bf",x"6e"),
  2364 => (x"ff",x"4b",x"87",x"c5"),
  2365 => (x"c1",x"0f",x"73",x"49"),
  2366 => (x"c4",x"49",x"75",x"7e"),
  2367 => (x"ce",x"c0",x"05",x"99"),
  2368 => (x"49",x"f2",x"c3",x"87"),
  2369 => (x"70",x"87",x"e4",x"e3"),
  2370 => (x"02",x"99",x"c2",x"49"),
  2371 => (x"c2",x"87",x"eb",x"c0"),
  2372 => (x"7e",x"bf",x"e4",x"f7"),
  2373 => (x"b7",x"c7",x"48",x"6e"),
  2374 => (x"cb",x"c0",x"03",x"a8"),
  2375 => (x"c1",x"48",x"6e",x"87"),
  2376 => (x"e8",x"f7",x"c2",x"80"),
  2377 => (x"87",x"d0",x"c0",x"58"),
  2378 => (x"c1",x"4a",x"66",x"c4"),
  2379 => (x"02",x"6a",x"82",x"e0"),
  2380 => (x"4b",x"87",x"c5",x"c0"),
  2381 => (x"0f",x"73",x"49",x"fe"),
  2382 => (x"fd",x"c3",x"7e",x"c1"),
  2383 => (x"87",x"eb",x"e2",x"49"),
  2384 => (x"99",x"c2",x"49",x"70"),
  2385 => (x"87",x"e6",x"c0",x"02"),
  2386 => (x"bf",x"e4",x"f7",x"c2"),
  2387 => (x"87",x"c9",x"c0",x"02"),
  2388 => (x"48",x"e4",x"f7",x"c2"),
  2389 => (x"d3",x"c0",x"78",x"c0"),
  2390 => (x"48",x"66",x"c4",x"87"),
  2391 => (x"70",x"80",x"e0",x"c1"),
  2392 => (x"02",x"bf",x"6e",x"7e"),
  2393 => (x"4b",x"87",x"c5",x"c0"),
  2394 => (x"0f",x"73",x"49",x"fd"),
  2395 => (x"fa",x"c3",x"7e",x"c1"),
  2396 => (x"87",x"f7",x"e1",x"49"),
  2397 => (x"99",x"c2",x"49",x"70"),
  2398 => (x"87",x"ea",x"c0",x"02"),
  2399 => (x"bf",x"e4",x"f7",x"c2"),
  2400 => (x"a8",x"b7",x"c7",x"48"),
  2401 => (x"87",x"c9",x"c0",x"03"),
  2402 => (x"48",x"e4",x"f7",x"c2"),
  2403 => (x"d3",x"c0",x"78",x"c7"),
  2404 => (x"48",x"66",x"c4",x"87"),
  2405 => (x"70",x"80",x"e0",x"c1"),
  2406 => (x"02",x"bf",x"6e",x"7e"),
  2407 => (x"4b",x"87",x"c5",x"c0"),
  2408 => (x"0f",x"73",x"49",x"fc"),
  2409 => (x"48",x"75",x"7e",x"c1"),
  2410 => (x"cc",x"98",x"f0",x"c3"),
  2411 => (x"98",x"70",x"58",x"a6"),
  2412 => (x"87",x"ce",x"c0",x"05"),
  2413 => (x"e0",x"49",x"da",x"c1"),
  2414 => (x"49",x"70",x"87",x"f1"),
  2415 => (x"c1",x"02",x"99",x"c2"),
  2416 => (x"e8",x"cf",x"87",x"f9"),
  2417 => (x"87",x"d0",x"c3",x"49"),
  2418 => (x"f7",x"c2",x"4b",x"70"),
  2419 => (x"50",x"c0",x"48",x"dc"),
  2420 => (x"97",x"dc",x"f7",x"c2"),
  2421 => (x"d2",x"c1",x"05",x"bf"),
  2422 => (x"05",x"66",x"c8",x"87"),
  2423 => (x"c1",x"87",x"cc",x"c0"),
  2424 => (x"c6",x"e0",x"49",x"da"),
  2425 => (x"02",x"98",x"70",x"87"),
  2426 => (x"e8",x"87",x"c0",x"c1"),
  2427 => (x"c3",x"49",x"4d",x"bf"),
  2428 => (x"b7",x"c8",x"99",x"ff"),
  2429 => (x"ff",x"b5",x"71",x"2d"),
  2430 => (x"73",x"87",x"f3",x"da"),
  2431 => (x"87",x"e4",x"c2",x"49"),
  2432 => (x"c0",x"02",x"98",x"70"),
  2433 => (x"f7",x"c2",x"87",x"c6"),
  2434 => (x"50",x"c1",x"48",x"dc"),
  2435 => (x"97",x"dc",x"f7",x"c2"),
  2436 => (x"d6",x"c0",x"05",x"bf"),
  2437 => (x"c3",x"49",x"75",x"87"),
  2438 => (x"ff",x"05",x"99",x"f0"),
  2439 => (x"da",x"c1",x"87",x"cd"),
  2440 => (x"c6",x"df",x"ff",x"49"),
  2441 => (x"05",x"98",x"70",x"87"),
  2442 => (x"c2",x"87",x"c0",x"ff"),
  2443 => (x"49",x"bf",x"e4",x"f7"),
  2444 => (x"c4",x"93",x"cc",x"4b"),
  2445 => (x"4b",x"6b",x"83",x"66"),
  2446 => (x"74",x"0f",x"73",x"71"),
  2447 => (x"e9",x"c0",x"02",x"9c"),
  2448 => (x"c0",x"02",x"6c",x"87"),
  2449 => (x"49",x"6c",x"87",x"e4"),
  2450 => (x"87",x"df",x"de",x"ff"),
  2451 => (x"99",x"c1",x"49",x"70"),
  2452 => (x"87",x"cb",x"c0",x"02"),
  2453 => (x"c2",x"4b",x"a4",x"c4"),
  2454 => (x"49",x"bf",x"e4",x"f7"),
  2455 => (x"c8",x"0f",x"4b",x"6b"),
  2456 => (x"c5",x"c0",x"02",x"84"),
  2457 => (x"ff",x"05",x"6c",x"87"),
  2458 => (x"02",x"6e",x"87",x"dc"),
  2459 => (x"c2",x"87",x"c8",x"c0"),
  2460 => (x"49",x"bf",x"e4",x"f7"),
  2461 => (x"f4",x"87",x"e9",x"f1"),
  2462 => (x"26",x"4d",x"26",x"8e"),
  2463 => (x"26",x"4b",x"26",x"4c"),
  2464 => (x"00",x"00",x"00",x"4f"),
  2465 => (x"00",x"00",x"00",x"10"),
  2466 => (x"00",x"00",x"00",x"00"),
  2467 => (x"00",x"00",x"00",x"00"),
  2468 => (x"00",x"00",x"00",x"00"),
  2469 => (x"00",x"00",x"00",x"00"),
  2470 => (x"ff",x"4a",x"71",x"1e"),
  2471 => (x"72",x"49",x"bf",x"c8"),
  2472 => (x"4f",x"26",x"48",x"a1"),
  2473 => (x"bf",x"c8",x"ff",x"1e"),
  2474 => (x"c0",x"c0",x"fe",x"89"),
  2475 => (x"a9",x"c0",x"c0",x"c0"),
  2476 => (x"c0",x"87",x"c4",x"01"),
  2477 => (x"c1",x"87",x"c2",x"4a"),
  2478 => (x"26",x"48",x"72",x"4a"),
  2479 => (x"5b",x"5e",x"0e",x"4f"),
  2480 => (x"71",x"0e",x"5d",x"5c"),
  2481 => (x"4c",x"d4",x"ff",x"4b"),
  2482 => (x"c0",x"48",x"66",x"d0"),
  2483 => (x"ff",x"49",x"d6",x"78"),
  2484 => (x"c3",x"87",x"d5",x"dd"),
  2485 => (x"49",x"6c",x"7c",x"ff"),
  2486 => (x"71",x"99",x"ff",x"c3"),
  2487 => (x"f0",x"c3",x"49",x"4d"),
  2488 => (x"a9",x"e0",x"c1",x"99"),
  2489 => (x"c3",x"87",x"cb",x"05"),
  2490 => (x"48",x"6c",x"7c",x"ff"),
  2491 => (x"66",x"d0",x"98",x"c3"),
  2492 => (x"ff",x"c3",x"78",x"08"),
  2493 => (x"49",x"4a",x"6c",x"7c"),
  2494 => (x"ff",x"c3",x"31",x"c8"),
  2495 => (x"71",x"4a",x"6c",x"7c"),
  2496 => (x"c8",x"49",x"72",x"b2"),
  2497 => (x"7c",x"ff",x"c3",x"31"),
  2498 => (x"b2",x"71",x"4a",x"6c"),
  2499 => (x"31",x"c8",x"49",x"72"),
  2500 => (x"6c",x"7c",x"ff",x"c3"),
  2501 => (x"ff",x"b2",x"71",x"4a"),
  2502 => (x"e0",x"c0",x"48",x"d0"),
  2503 => (x"02",x"9b",x"73",x"78"),
  2504 => (x"7b",x"72",x"87",x"c2"),
  2505 => (x"4d",x"26",x"48",x"75"),
  2506 => (x"4b",x"26",x"4c",x"26"),
  2507 => (x"26",x"1e",x"4f",x"26"),
  2508 => (x"5b",x"5e",x"0e",x"4f"),
  2509 => (x"86",x"f8",x"0e",x"5c"),
  2510 => (x"a6",x"c8",x"1e",x"76"),
  2511 => (x"87",x"fd",x"fd",x"49"),
  2512 => (x"4b",x"70",x"86",x"c4"),
  2513 => (x"a8",x"c4",x"48",x"6e"),
  2514 => (x"87",x"fb",x"c2",x"03"),
  2515 => (x"f0",x"c3",x"4a",x"73"),
  2516 => (x"aa",x"d0",x"c1",x"9a"),
  2517 => (x"c1",x"87",x"c7",x"02"),
  2518 => (x"c2",x"05",x"aa",x"e0"),
  2519 => (x"49",x"73",x"87",x"e9"),
  2520 => (x"c3",x"02",x"99",x"c8"),
  2521 => (x"87",x"c6",x"ff",x"87"),
  2522 => (x"9c",x"c3",x"4c",x"73"),
  2523 => (x"c1",x"05",x"ac",x"c2"),
  2524 => (x"66",x"c4",x"87",x"c4"),
  2525 => (x"71",x"31",x"c9",x"49"),
  2526 => (x"4a",x"66",x"c4",x"1e"),
  2527 => (x"c2",x"92",x"cc",x"c1"),
  2528 => (x"72",x"49",x"ec",x"f7"),
  2529 => (x"c1",x"cd",x"fe",x"81"),
  2530 => (x"ff",x"49",x"d8",x"87"),
  2531 => (x"c8",x"87",x"d9",x"da"),
  2532 => (x"e4",x"c2",x"1e",x"c0"),
  2533 => (x"e6",x"fd",x"49",x"e4"),
  2534 => (x"d0",x"ff",x"87",x"d9"),
  2535 => (x"78",x"e0",x"c0",x"48"),
  2536 => (x"1e",x"e4",x"e4",x"c2"),
  2537 => (x"c1",x"4a",x"66",x"cc"),
  2538 => (x"f7",x"c2",x"92",x"cc"),
  2539 => (x"81",x"72",x"49",x"ec"),
  2540 => (x"87",x"d7",x"cb",x"fe"),
  2541 => (x"ac",x"c1",x"86",x"cc"),
  2542 => (x"87",x"cb",x"c1",x"05"),
  2543 => (x"fd",x"49",x"ee",x"c0"),
  2544 => (x"c4",x"87",x"c9",x"e3"),
  2545 => (x"31",x"c9",x"49",x"66"),
  2546 => (x"66",x"c4",x"1e",x"71"),
  2547 => (x"92",x"cc",x"c1",x"4a"),
  2548 => (x"49",x"ec",x"f7",x"c2"),
  2549 => (x"cb",x"fe",x"81",x"72"),
  2550 => (x"e4",x"c2",x"87",x"f0"),
  2551 => (x"66",x"c8",x"1e",x"e4"),
  2552 => (x"92",x"cc",x"c1",x"4a"),
  2553 => (x"49",x"ec",x"f7",x"c2"),
  2554 => (x"c9",x"fe",x"81",x"72"),
  2555 => (x"49",x"d7",x"87",x"de"),
  2556 => (x"87",x"f4",x"d8",x"ff"),
  2557 => (x"c2",x"1e",x"c0",x"c8"),
  2558 => (x"fd",x"49",x"e4",x"e4"),
  2559 => (x"cc",x"87",x"d1",x"e4"),
  2560 => (x"48",x"d0",x"ff",x"86"),
  2561 => (x"f8",x"78",x"e0",x"c0"),
  2562 => (x"26",x"4c",x"26",x"8e"),
  2563 => (x"1e",x"4f",x"26",x"4b"),
  2564 => (x"b7",x"c4",x"4a",x"71"),
  2565 => (x"87",x"ce",x"03",x"aa"),
  2566 => (x"cc",x"c1",x"49",x"72"),
  2567 => (x"ec",x"f7",x"c2",x"91"),
  2568 => (x"81",x"c8",x"c1",x"81"),
  2569 => (x"4f",x"26",x"79",x"c0"),
  2570 => (x"5c",x"5b",x"5e",x"0e"),
  2571 => (x"86",x"fc",x"0e",x"5d"),
  2572 => (x"d4",x"ff",x"4a",x"71"),
  2573 => (x"d4",x"4c",x"c0",x"4b"),
  2574 => (x"b7",x"c3",x"4d",x"66"),
  2575 => (x"c2",x"c2",x"01",x"ad"),
  2576 => (x"02",x"9a",x"72",x"87"),
  2577 => (x"1e",x"87",x"ec",x"c0"),
  2578 => (x"cc",x"c1",x"49",x"75"),
  2579 => (x"ec",x"f7",x"c2",x"91"),
  2580 => (x"c8",x"80",x"71",x"48"),
  2581 => (x"66",x"c4",x"58",x"a6"),
  2582 => (x"fb",x"c2",x"fe",x"49"),
  2583 => (x"70",x"86",x"c4",x"87"),
  2584 => (x"87",x"d4",x"02",x"98"),
  2585 => (x"c8",x"c1",x"49",x"6e"),
  2586 => (x"6e",x"79",x"c1",x"81"),
  2587 => (x"69",x"81",x"c8",x"49"),
  2588 => (x"75",x"87",x"c5",x"4c"),
  2589 => (x"87",x"d7",x"fe",x"49"),
  2590 => (x"c8",x"48",x"d0",x"ff"),
  2591 => (x"7b",x"dd",x"78",x"e1"),
  2592 => (x"ff",x"c3",x"48",x"74"),
  2593 => (x"74",x"7b",x"70",x"98"),
  2594 => (x"29",x"b7",x"c8",x"49"),
  2595 => (x"ff",x"c3",x"48",x"71"),
  2596 => (x"74",x"7b",x"70",x"98"),
  2597 => (x"29",x"b7",x"d0",x"49"),
  2598 => (x"ff",x"c3",x"48",x"71"),
  2599 => (x"74",x"7b",x"70",x"98"),
  2600 => (x"28",x"b7",x"d8",x"48"),
  2601 => (x"7b",x"c0",x"7b",x"70"),
  2602 => (x"7b",x"7b",x"7b",x"7b"),
  2603 => (x"7b",x"7b",x"7b",x"7b"),
  2604 => (x"ff",x"7b",x"7b",x"7b"),
  2605 => (x"e0",x"c0",x"48",x"d0"),
  2606 => (x"dc",x"1e",x"75",x"78"),
  2607 => (x"cc",x"d6",x"ff",x"49"),
  2608 => (x"fc",x"86",x"c4",x"87"),
  2609 => (x"26",x"4d",x"26",x"8e"),
  2610 => (x"26",x"4b",x"26",x"4c"),
  2611 => (x"00",x"00",x"00",x"4f"),
  2612 => (x"ff",x"ff",x"ff",x"ff"),
  2613 => (x"ff",x"ff",x"ff",x"ff"),
  2614 => (x"ff",x"ff",x"ff",x"ff"),
  2615 => (x"ff",x"ff",x"ff",x"ff"),
  2616 => (x"00",x"00",x"28",x"e4"),
  2617 => (x"33",x"49",x"56",x"53"),
  2618 => (x"20",x"20",x"38",x"32"),
  2619 => (x"00",x"4d",x"4f",x"52"),
  2620 => (x"00",x"00",x"1b",x"d3"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

